���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.6.1�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy._core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��	RestingBP��Cholesterol��	FastingBS��MaxHR��ExerciseAngina��Oldpeak��ChestPainType_ASY��ChestPainType_ATA��ChestPainType_NAP��ChestPainType_TA��RestingECG_LVH��RestingECG_Normal��RestingECG_ST��ST_Slope_Down��ST_Slope_Flat��ST_Slope_Up�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��h3�f8�����R�(KhXNNNJ����J����K t�b�C              �?�t�bh\h'�scalar���hWC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hK�
node_count�K�nodes�h)h,K ��h.��R�(KKᅔh3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h�hWK ��h�hWK��h�hWK��h�hiK��h�hiK ��h�hWK(��h�hiK0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@8         h                    �?j8je3�?�           ��@                                   �?�6tT�.�?�            �u@                                   @M@j�'�=z�?%            �P@                                  �^@|��?���?             ;@               
                   Pm@      �?             (@                                 �`@ףp=
�?             $@       ������������������������       �                     @               	                   �W@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                  �b@������?	             .@                                 �]@d}h���?             ,@                                ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?                                   @P@$�q-�?            �C@       ������������������������       �                     ;@                                   �P@      �?             (@        ������������������������       �                      @                                  �q@ףp=
�?             $@       ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               Y                    �?Df/��?�            �q@              X                 ���@ wVX(6�?�            `n@              W                   �g@T(y2��?�            �m@              H                 ����?86��Z�?�            �m@               5                   `_@�]��?�            �i@        !       2                    _@����!p�?:             V@       "       )                 833�?P��BNֱ?6            �T@       #       (       	             �?�}��L�?0            �R@       $       %                   pc@������?             B@       ������������������������       �                     5@        &       '                   �c@��S�ۿ?	             .@        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                    �C@        *       /                    �?      �?              @       +       ,                   @\@      �?             @        ������������������������       �                     �?        -       .                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        0       1                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        3       4                    �K@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        6       G                    �?���<_�?M            �]@       7       B                   �b@Pa�	�?B            �X@       8       9                   �c@p�C��?;            �V@       ������������������������       �        %             M@        :       ;                   �c@�FVQ&�?            �@@        ������������������������       �                     �?        <       =                    @I@      �?             @@       ������������������������       �                     9@        >       A       
             �?؇���X�?             @        ?       @                     J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        C       F                    m@      �?              @        D       E                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        I       P                    �L@��a�n`�?             ?@       J       K                    �?�����?             5@       ������������������������       �                     1@        L       O                    �?      �?             @       M       N                   pe@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        Q       T                    �?      �?             $@       R       S                   �k@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        U       V                 `ff�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Z       g       	             �?��
ц��?            �C@       [       f                    �?���Q��?             >@       \       ]                    �?X�Cc�?             <@        ������������������������       �                     @        ^       e                   Pd@ �o_��?             9@       _       `                    @M@ףp=
�?             4@        ������������������������       �                      @        a       b                   `_@r�q��?	             (@        ������������������������       �                     @        c       d                 ����?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        i       �                   �b@��SA_�?�             x@       j       �                    �?l{��b��?�            �s@       k       �                    �?���>4��?�             l@        l       �                 ����?�?�'�@�?5             S@       m       �                    �O@z�G�z�?             D@       n       q                    @G@     ��?             @@        o       p                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        r       w                   `X@@4և���?             <@        s       t                    �?�q�q�?             @        ������������������������       �                     �?        u       v                   @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       y                    �M@`2U0*��?             9@       ������������������������       �                     ,@        z       {       
             �?�C��2(�?             &@       ������������������������       �                      @        |                           �?�q�q�?             @       }       ~                   ``@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�X�<ݺ?             B@       �       �                    �?�C��2(�?             6@        ������������������������       �                      @        �       �                    �?؇���X�?	             ,@        ������������������������       �                      @        �       �                   �Z@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �        	             ,@        �       �                    �?����?Y            �b@        �       �                    �?�㙢�c�?             7@        �       �                    �?���|���?             &@        ������������������������       �                     @        �       �                   �q@      �?              @       �       �                 `ff�?�q�q�?             @       �       �       	             �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �l@0{�v��?I            @_@       �       �                 ����?L������?(            @R@        ������������������������       �                     8@        �       �                   @l@ZՏ�m|�?            �H@       �       �                   �g@�q��/��?             G@        ������������������������       �                     5@        �       �                 ����?z�G�z�?             9@        �       �                    �K@      �?             $@        ������������������������       �                     @        �       �                   �a@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     @        �       �                    �? pƵHP�?!             J@        ������������������������       �                     $@        �       �                    @I@�Ń��̧?             E@        �       �                    �?      �?              @        �       �                   @`@      �?             @       �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     A@        �       �                   �`@�����?5             W@       ������������������������       �        ,             S@        �       �                    n@      �?	             0@       ������������������������       �                     $@        �       �                   pa@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�Cc�?+            �Q@       �       �                    �?��+��?            �B@        �       �                     H@�t����?             1@       �       �                 ����?ףp=
�?             $@        ������������������������       �                     @        �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `]@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �L@�z�G��?             4@       ������������������������       �                     "@        �       �                   �c@�eP*L��?             &@        ������������������������       �                     @        �       �                 033�?؇���X�?             @        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `q@"pc�
�?            �@@       �       �                   c@����X�?             5@        ������������������������       �                      @        �       �                    q@���y4F�?             3@       �       �                    �?      �?
             0@       �       �                    �?"pc�
�?             &@       �       �                    @H@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �t�b�values�h)h,K ��h.��R�(KK�KK��hi�B  ���Y��?t�S��?[�~�u��?J��/�?|��|�?�|���?{	�%���?	�%����?      �?      �?�������?�������?              �?�������?�������?      �?                      �?      �?        wwwwww�?�?I�$I�$�?۶m۶m�?�������?333333�?      �?                      �?      �?                      �?;�;��?�؉�؉�?              �?      �?      �?      �?        �������?�������?              �?      �?      �?              �?      �?        � &W��?G}g����?k~X�<�?�<ݚ�?�F��F��?�5�5�?�Z܄��?h *�3�?p�14���?��,�?/�袋.�?]t�E�?��FS���?���ˊ��?�_,�Œ�?O贁N�?�q�q�?�q�q�?      �?        �������?�?              �?      �?              �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        333333�?�������?      �?                      �?+����/�?��/���?|���?|���?��K��K�?h�h��?      �?        >����?|���?              �?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?      �?      �?      �?      �?                      �?      �?              �?        �c�1��?�s�9��?=��<���?�a�a�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?�������?�������?              �?      �?        �������?�������?              �?      �?                      �?              �?�;�;�?�؉�؉�?�������?333333�?�m۶m��?%I�$I��?      �?        �Q����?
ףp=
�?�������?�������?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?        0���?�?�H	9��?�&��jq�?${�ґ�?�$I�$I�?n۶m۶�?y�5���?������?�������?�������?      �?      �?      �?      �?      �?                      �?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        {�G�z�?���Q��?              �?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        �q�q�?��8��8�?F]t�E�?]t�E�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?              �?�g�`�|�?S�n0�?d!Y�B�?�7��Mo�?F]t�E�?]t�E]�?              �?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?                      �?;�O��n�?V-��?����?�Ǐ?~�?              �?9/����?�>4և��?��Mozӻ?�B����?              �?�������?�������?      �?      �?              �?�������?UUUUUU�?      �?                      �?              �?      �?        ;�;��?'vb'vb�?              �?�a�a�?��<��<�?      �?      �?      �?      �?      �?      �?              �?      �?                      �?              �?              �?d!Y�B�?zӛ����?              �?      �?      �?              �?UUUUUU�?�������?      �?                      �?�m۶m��?%I�$I��?�S�n�?*�Y7�"�?�������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        ffffff�?333333�?      �?        ]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?F]t�E�?/�袋.�?�$I�$I�?�m۶m��?      �?        (������?6��P^C�?      �?      �?F]t�E�?/�袋.�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKᅔh��B@8         b                    �?4�5����?�           ��@               +                    �?R�чf��?�            �u@                                  @L@��t��?�            �l@                                  �?�8���?k            �e@                                  @h�����?f             e@              	       
             �? Df@��?e            �d@                                 �g@` A�c̭?>             Y@       ������������������������       �        =            @X@        ������������������������       �                     @        
                          �m@����e��?'            �P@       ������������������������       �                     F@                                   �?���7�?             6@        ������������������������       �                     &@                                   �?�C��2(�?             &@                                 �c@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                   �G@      �?             @        ������������������������       �                      @                                   �?      �?             @        ������������������������       �                     �?                                  e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               (                 `ff�?>4և���?              L@              %                   ht@R���Q�?             D@              "                   �?��G���?            �B@              !                    �? �Cc}�?             <@                                   �c@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �        	             0@        #       $                    �M@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        &       '                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        )       *                    �?      �?	             0@        ������������������������       �                      @        ������������������������       �                     ,@        ,       O                    �?"� ���?O            @]@       -       H                    �?v�X��?<             V@       .       G                 ��� @:���W�?*            �M@       /       4                   �h@��V�I��?"            �G@        0       3                    �?�IєX�?             1@        1       2                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             *@        5       <                   �_@�q�q�?             >@        6       ;                     N@�<ݚ�?             "@        7       8                    �L@�q�q�?             @        ������������������������       �                     �?        9       :                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        =       >                    �?؇���X�?             5@        ������������������������       �                     "@        ?       @                   m@      �?             (@        ������������������������       �                     @        A       B                   Pa@      �?             @        ������������������������       �                      @        C       F       	             �?      �?             @       D       E                    @E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        I       N                   c@д>��C�?             =@       J       M                    �?`2U0*��?             9@        K       L                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     @        P       Q                    �?8^s]e�?             =@        ������������������������       �                     "@        R       Y       
             �?�G�z��?             4@        S       T                 ����?���!pc�?             &@        ������������������������       �                     �?        U       V                   �c@z�G�z�?             $@       ������������������������       �                     @        W       X                   �b@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        Z       _                    �?�q�q�?             "@       [       ^                    @�q�q�?             @       \       ]                   pc@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        `       a                    ^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        c       �                    �?�#�k���?�            0x@        d       �                 ����?X�Emq�?b            �c@        e       |                    �?��i#[�?0             U@       f       s                    �?<ݚ�?(             R@       g       l                    �?�:�]��?            �I@       h       i                   �k@`���i��?             F@       ������������������������       �                     =@        j       k                   �l@��S�ۿ?	             .@        ������������������������       �                     �?        ������������������������       �                     ,@        m       r                   �c@և���X�?             @       n       o                    �?z�G�z�?             @        ������������������������       �                     @        p       q                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        t       {                 ����?�ՙ/�?	             5@       u       z                   �f@X�<ݚ�?             2@       v       y                    p@�θ�?             *@        w       x                    @H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        }       �                    �?      �?             (@       ~                           �E@�q�q�?             "@        ������������������������       �                      @        �       �                   ``@և���X�?             @       �       �                 ,33ӿz�G�z�?             @        ������������������������       �                      @        �       �                   `@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���?2            �R@       �       �                   �U@�j��b�?'            �M@        ������������������������       �                     �?        �       �                    �R@��ϭ�*�?&             M@       �       �                   ``@l�b�G��?%            �L@       �       �                 ����?г�wY;�?             A@        �       �                    �?z�G�z�?             @       �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     =@        �       �                    x@�LQ�1	�?             7@       �       �                    �?�C��2(�?             6@        �       �                    �O@      �?              @       �       �                   �k@؇���X�?             @        ������������������������       �                     @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?     ��?             0@       �       �                   �_@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �r@�q�q�?             @       �       �                   �a@      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?x�}b~|�?�            �l@       �       �                   `_@�$�����?g            @d@       �       �                    �?��S�ۿ?;            �V@       �       �                    �?�L���?3            �R@        ������������������������       �                     $@        �       �                    �H@     ��?,             P@        ������������������������       �        	             *@        �       �                   xt@�t����?#            �I@       �       �                   `l@dP-���?!            �G@        ������������������������       �                     1@        �       �                    �?�r����?             >@        �       �                    �?      �?              @        �       �                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `\@r�q��?             @        �       �                   @X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `m@�C��2(�?             6@        ������������������������       �                     �?        �       �                    �O@���N8�?             5@       ������������������������       �        
             4@        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        �       �                    �?tk~X��?,             R@       �       �                   0i@`��:�?%            �N@        �       �                   �b@     ��?
             0@        ������������������������       �                     @        �       �                 ����?�q�q�?             (@        ������������������������       �                      @        �       �                    �I@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                   pc@�����H�?            �F@       �       �                   �l@�}�+r��?             C@        �       �                   �k@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     <@        �       �                   xu@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   Pm@"pc�
�?             &@       ������������������������       �                      @        �       �                    @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        &            �P@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B   Np	�?���Gw{�?ٮ�n^��?N��"C��?�_�T>��?�����?j��FX�?a���{�?�m۶m��?�$I�$I�?c��7�:�?��k���?
ףp=
�?���Q��?      �?                      �?�>����?|���?      �?        �.�袋�?F]t�E�?      �?        ]t�E�?F]t�E�?�q�q�?�q�q�?              �?      �?              �?                      �?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?�������?�������?#�u�)��?v�)�Y7�?%I�$I��?۶m۶m�?      �?      �?      �?                      �?      �?        r�q��?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?��)��)�?�6k�6k�?颋.���?�.�袋�?A�Iݗ��?_[4��?r1����?G}g����?�?�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?|a���?a���{�?{�G�z�?���Q��?      �?      �?      �?                      �?              �?      �?        |a���?	�=����?      �?        �������?�������?F]t�E�?t�E]t�?              �?�������?�������?      �?        333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        \���o�?)��:��?�}�	��?5�x+��?�a�a�?�<��<��?�q�q�?��8��8�?}}}}}}�?�?F]t�E�?F]t�E�?      �?        �������?�?              �?      �?        �$I�$I�?۶m۶m�?�������?�������?      �?              �?      �?      �?                      �?              �?�a�a�?�<��<��?�q�q�?r�q��?�؉�؉�?ى�؉��?      �?      �?              �?      �?                      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?ƒ_,���?O贁N�?��/���?�N��?      �?        |a���?����=�?p�}��?�Gp��?�?�?�������?�������?      �?      �?              �?      �?                      �?              �?Y�B��?��Moz��?F]t�E�?]t�E�?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?              �?      �?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?Lg1��t�?�YLg1�?X�<ݚ�?uk~X��?�?�������?L�Ϻ��?}���g�?              �?      �?      �?              �?�?<<<<<<�?W�+�ɵ?�����F�?              �?�?�������?      �?      �?      �?      �?              �?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?F]t�E�?]t�E�?      �?        �a�a�?��y��y�?              �?      �?              �?      �?              �?      �?                      �?9��8���?r�q��?XG��).�?*.�u��?      �?      �?              �?�������?�������?              �?ffffff�?333333�?              �?      �?        �q�q�?�q�q�?(�����?�5��P�?�������?�������?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?        F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�/         V                    �?p�Vv���?�           ��@                                  �O@¦	^_�?�            Pu@                                   �?������?             >@                                  �?`�Q��?             9@                     	             �?��S���?             .@                                  �?���|���?             &@                                433�?և���X�?             @        ������������������������       �                     @        	       
                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?ףp=
�?             $@        ������������������������       �                     @                                `ff@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               C                    �?Z�WUL��?�            ps@               "                    �?C7�J�?G            �[@                                   �?      �?             8@        ������������������������       �                     @                                   [@R���Q�?             4@        ������������������������       �                     �?               !                 ����?�KM�]�?             3@                                ����?"pc�
�?             &@                                 �q@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        #       4                 ����?RB)��.�?8            �U@        $       %                   pk@#z�i��?            �D@        ������������������������       �                     &@        &       -                    �?��S���?             >@       '       (                 ����?�q�q�?             2@        ������������������������       �                     "@        )       ,                    �L@�q�q�?             "@        *       +                     E@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        .       /                   �]@�q�q�?             (@        ������������������������       �                     @        0       3                    �?      �?              @       1       2                   �q@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        5       B                   �`@�:�^���?            �F@        6       A                    `@�q�q�?             (@       7       8                    �?z�G�z�?
             $@        ������������������������       �                     @        9       <       
             �?����X�?             @       :       ;                    @I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        =       >                    �?�q�q�?             @        ������������������������       �                     �?        ?       @                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �@@        D       U                    @0�,���?~             i@       E       T                   �g@�ʱ�O+�?|            �h@       F       G                   �?����e��?{            �h@       ������������������������       �        f            �d@        H       S                   a@��a�n`�?             ?@       I       R       
             �?r�q��?             2@       J       M                   �a@d}h���?	             ,@        K       L                   pa@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        N       Q                    j@�����H�?             "@        O       P       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             *@        ������������������������       �                     �?        ������������������������       �                      @        W       �                    �?�x�V�"�?           �x@        X       _                   �_@v�(��O�?a            �b@        Y       ^                   �^@P�Lt�<�?             C@        Z       [                 033�?�}�+r��?             3@       ������������������������       �        	             .@        \       ]                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        `       y                   �a@     ��?F             \@       a       l                    �?<�\`*��?5             U@       b       i                    �?     ��?(             P@       c       h                    �?P���Q�?             D@       d       e                 hff�?@4և���?             <@       ������������������������       �                     9@        f       g                   pe@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        j       k                    @L@�q�q�?             8@       ������������������������       �                     0@        ������������������������       �                      @        m       v                 ����?�G�z��?             4@       n       o                   �\@�n_Y�K�?             *@        ������������������������       �                     @        p       u                    �?����X�?             @       q       r                     G@      �?             @        ������������������������       �                     �?        s       t                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        w       x                   `v@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        z       �                    �?����X�?             <@       {       |                    �?��2(&�?             6@       ������������������������       �                     *@        }       �                    �O@�q�q�?             "@       ~       �                   �b@؇���X�?             @               �                    l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?r�q��?             @       �       �                    @P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�>����?�            `n@        �       �                   Pd@�[|x��?*            �O@       �       �                   P`@�.ߴ#�?(            �N@       ������������������������       �                     E@        �       �                   �b@�S����?             3@       ������������������������       �        	             .@        �       �                 ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0c@0��Q'�?w            �f@       �       �                   i@���1j	�?r            �e@        ������������������������       �        $             M@        �       �                    j@x�}b~|�?N            �\@        �       �                   �i@      �?              @       �       �                     L@      �?             @        ������������������������       �                      @        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����?H            �Z@       �       �                    \@(;L]n�?%             N@        �       �                    �J@�C��2(�?
             &@        �       �                    Z@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?@�E�x�?            �H@       �       �                    �?XB���?             =@        ������������������������       �                     @        �       �                     H@`2U0*��?             9@        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     4@        �       �                    @I@���.�6�?#             G@        �       �                    �H@؇���X�?
             ,@       �       �                   �_@$�q-�?	             *@       ������������������������       �                     @        �       �                   �m@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    `@      �?             @@        �       �                    @O@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �m@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  w
��,@�?�z�����?��Zk���?�RJ)���?�?wwwwww�?{�G�z�?��(\���?�������?�?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?                      �?�������?�������?              �?�������?�������?              �?      �?                      �?h��p��?a��<���?��k߰�?�yJ���?      �?      �?      �?        333333�?333333�?              �?�k(���?(�����?/�袋.�?F]t�E�?�������?�������?      �?                      �?              �?      �?        ���)k��?S֔5eM�?ە�]���?�+Q��?              �?�������?�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?l�l��?}�'}�'�?UUUUUU�?UUUUUU�?�������?�������?              �?�$I�$I�?�m۶m��?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?Ez�rv�?g��1��?}i�0V[�?gв�9��?�>����?|���?      �?        �s�9��?�c�1Ƹ?�������?UUUUUU�?I�$I�$�?۶m۶m�?333333�?�������?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?              �?                      �?              �?�����?�y�L�R�?O贁N�?Y�%�X�?(�����?���k(�?(�����?�5��P�?              �?      �?      �?      �?                      �?              �?      �?      �?=��<���?�a�a�?      �?      �?ffffff�?�������?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?�m۶m��?t�E]t�?��.���?              �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        h/�����?�Kh/��?EQEQ�?]�u]�u�?XG��).�?�K�`m�?              �?^Cy�5�?(������?              �?      �?      �?      �?                      �?      �?        �'}�'}�?[�[��?qG�wĭ?�;⎸#�?              �?Lg1��t�?�YLg1�?      �?      �?      �?      �?              �?      �?      �?              �?      �?              �?        �V�9�&�?��`��}�?�?�������?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?9/���?և���X�?�{a���?GX�i���?              �?{�G�z�?���Q��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?Y�B��?���7���?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?              �?UUUUUU�?�������?      �?                      �?      �?              �?      �?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?      �?              �?333333�?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKᅔh��B@8         t                    �?U�ք�?�           ��@               ?                 pff�?:"Z��?�            �u@              8                    �?���B���?�            @p@                                  �?��[�\�?�             n@              
                    �?P�Lt�<�?            �g@                                   �?��v$���?)            �N@       ������������������������       �        #             J@               	                   P`@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                  �g@0Ƭ!sĮ?V             `@                                 �t@     p�?U             `@                     
             �?������?T            �_@                                  �?����e��?/            �P@       ������������������������       �        ,            �O@                                  �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        %             N@        ������������������������       �                      @        ������������������������       �                     �?                                   �F@�q�q�?$            �I@        ������������������������       �                     @               3                    �?��Hg���?            �F@                                   �?�t����?             A@                                   �?���Q��?             $@                                 �q@�q�q�?             "@                                  @I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        !       &       
             �?r�q��?             8@        "       #                 ����?�q�q�?             @        ������������������������       �                     @        $       %                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        '       (                    �L@�����H�?             2@        ������������������������       �                     "@        )       0                    �?�<ݚ�?             "@       *       /                     N@؇���X�?             @        +       ,                   �]@�q�q�?             @        ������������������������       �                     �?        -       .                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        1       2                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       5                    �M@�C��2(�?             &@       ������������������������       �                     @        6       7                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        9       >                 ����?D�n�3�?             3@       :       ;                    �?d}h���?	             ,@       ������������������������       �                     $@        <       =                   pb@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        @       i                    �?��>4և�?7             U@       A       T                 `ff�?�\����?+            �P@       B       S                   `b@ҳ�wY;�?             A@       C       D                   �c@և���X�?             <@        ������������������������       �                     @        E       R                    �?��H�}�?             9@       F       G                    �?�\��N��?             3@        ������������������������       �                     @        H       M                    �?����X�?             ,@        I       L                    �?      �?              @       J       K                   a@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        N       O       	             �?r�q��?             @       ������������������������       �                     @        P       Q                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        U       d                    �?     ��?             @@       V       a                    
@���B���?             :@       W       ^                   @a@r�q��?             8@       X       Y                   �g@      �?             0@       ������������������������       �                     "@        Z       ]                   �`@؇���X�?             @       [       \                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        _       `                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        b       c                 033@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       f       
             �?�q�q�?             @        ������������������������       �                      @        g       h                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        j       k                    �?�����H�?             2@        ������������������������       �                     @        l       m                   @_@"pc�
�?	             &@        ������������������������       �                     �?        n       s                    �?ףp=
�?             $@        o       p       
             �?�q�q�?             @        ������������������������       �                     �?        q       r                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        u       �                   �f@f�ȭ��?�            `x@       v       �                    �?�r���?�            �w@       w       �                    a@�,�bON�?�            0p@       x       }                    �?�Q��k�?j             d@        y       |                   �`@��S���?             .@       z       {                 ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                    �?(9jl8&�?_             b@               �                    �?     ��?             @@       �       �                   �_@�q�q�?             8@       �       �                    �?�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@        �       �                    �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?ЮN
��?G            @\@       �       �                   i@X'"7��?D             [@        ������������������������       �                     E@        �       �                    \@�U�=���?)            �P@        �       �                    @J@PN��T'�?             ;@        ������������������������       �                     *@        �       �                    �?����X�?
             ,@        �       �                    �?      �?             @        �       �                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@ףp=
�?             $@        �       �                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �_@ ���J��?            �C@       �       �                   �\@P���Q�?             4@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �        
             3@        �       �                   �Z@z�G�z�?             @       �       �                   b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �K@v�C��?A            �X@       �       �                   �b@���Q��?'            �K@        �       �                    �?z�G�z�?             9@        �       �                    �?$�q-�?             *@       ������������������������       �                     &@        �       �                    h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?             (@        ������������������������       �                     @        �       �                   `]@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �e@*;L]n�?             >@        ������������������������       �                      @        �       �                    �?��>4և�?             <@        �       �                 ����?ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    `@X�<ݚ�?             2@        �       �                    �E@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pf@�	j*D�?	             *@       �       �                 ����?      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?fP*L��?             F@        �       �                    �?�����?             3@        ������������������������       �                     $@        �       �                   �n@�q�q�?             "@       �       �                   Pc@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@`2U0*��?             9@        �       �                   `@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                    �?Hn�.P��?J             _@       �       �                    �?@3����?@             [@       ������������������������       �        3            @V@        �       �                   �o@�KM�]�?             3@       ������������������������       �                     0@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @\@      �?
             0@        �       �                     Q@z�G�z�?             @       �       �                    V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �t�b��,     h�h)h,K ��h.��R�(KK�KK��hi�B  ᓔ��?�5�;��?��)kʚ�?���)k��?��؉���?ى�؉��?�R��R��?�������?���k(�?(�����?.�u�y�?;ڼOqɐ?      �?        �q�q�?�q�q�?              �?      �?        ����?����?     @�?      �?�������?AA�?�>����?|���?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?UUUUUU�?UUUUUU�?      �?        ��I��I�?؂-؂-�?�������?�������?333333�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?�q�q�?9��8���?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?F]t�E�?]t�E�?              �?      �?      �?              �?      �?        (������?l(�����?۶m۶m�?I�$I�$�?              �?      �?      �?      �?                      �?      �?        I�$I�$�?۶m۶m�?>����?���>��?�������?�������?�$I�$I�?۶m۶m�?              �?{�G�z�?
ףp=
�?y�5���?�5��P�?              �?�m۶m��?�$I�$I�?      �?      �?�m۶m��?�$I�$I�?              �?      �?                      �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?              �?      �?ى�؉��?��؉���?UUUUUU�?�������?      �?      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �q�q�?�q�q�?              �?F]t�E�?/�袋.�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?ڞ�ٞ��?J��I���?>�˱
�?��S���?���O�?�}+�v��?�������?�������?�������?�?      �?      �?      �?                      �?              �?�[���?�Ő��?      �?      �?�������?UUUUUU�?(�����?�k(���?      �?                      �?333333�?�������?              �?      �?              �?        4��A�/�?m���M�?B{	�%��?Lh/����?              �?e�M6�d�?�M6�d��?h/�����?&���^B�?              �?�$I�$I�?�m۶m��?      �?      �?      �?      �?              �?      �?              �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�A�A�?��-��-�?�������?ffffff�?�������?�������?      �?                      �?              �?              �?�������?�������?      �?      �?              �?      �?                      �?1ogH���?gH���?333333�?�������?�������?�������?�؉�؉�?;�;��?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?�������?""""""�?      �?        I�$I�$�?۶m۶m�?�������?�������?              �?      �?        r�q��?�q�q�?�������?�������?      �?                      �?vb'vb'�?;�;��?      �?      �?      �?                      �?              �?]t�E]�?颋.���?^Cy�5�?Q^Cy��?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?{�G�z�?���Q��?�������?�������?              �?      �?                      �?�c�1ƨ?t�9�s�?h/�����?���Kh�?              �?(�����?�k(���?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B@>         �       	             �?4�5����?�           ��@              �                    �?�)��V�?�           ��@              B                    �?,g0M�h�?�            @x@               %                   �b@r�qG�?_             b@                                  �?H;T*St�?A            �X@               	                 ����?և���X�?
             ,@                                   ^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        
                           �?�z�G��?             $@                                 @_@�<ݚ�?             "@                                   �P@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                ����?�8��8��?7             U@        ������������������������       �                     A@                                    �?�:pΈ��?              I@                                 �[@�+$�jP�?             ;@        ������������������������       �                      @                                  �m@�d�����?             3@                               hff@�q�q�?	             .@                                  �?X�<ݚ�?             "@                                   �O@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �e@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        !       $                    �?���}<S�?             7@        "       #                    �M@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             2@        &       3                   a@\X��t�?             G@       '       ,                   �Q@�<ݚ�?             ;@        (       +                    �?z�G�z�?             @        )       *                   0d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        -       .                    @G@�C��2(�?             6@        ������������������������       �                     &@        /       0                   `\@"pc�
�?             &@        ������������������������       �                     �?        1       2                    e@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        4       =                    �?�d�����?             3@       5       6                   �a@�	j*D�?             *@        ������������������������       �                     @        7       :       
             �?և���X�?             @        8       9                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ;       <                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        >       A                 `ff�?r�q��?             @        ?       @                   pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        C       �                   �a@\#r��?�            �n@       D       E                   �Y@�H��?�?n             e@        ������������������������       �                     @        F       Y                    �G@؇���X�?i             d@        G       H                    �?$��m��?             :@        ������������������������       �                     @        I       P                    �?��+7��?             7@        J       K                   �`@և���X�?             @        ������������������������       �                     @        L       O                    �?      �?             @       M       N                   pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        Q       R                    �?     ��?             0@        ������������������������       �                     @        S       X                    �?�q�q�?             "@       T       W                    �?և���X�?             @       U       V                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        Z       [                    �?�Aʑ���?W            �`@        ������������������������       �        
             *@        \       s                   `\@Xny��?M            �^@        ]       ^                   �i@      �?             @@        ������������������������       �                     "@        _       j                   `[@�LQ�1	�?             7@       `       e                    �?������?
             1@       a       d                 433�?�8��8��?             (@        b       c                   `Y@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        f       g                    �?���Q��?             @        ������������������������       �                     �?        h       i                   (q@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        k       l                   �n@�q�q�?             @        ������������������������       �                      @        m       n                    �I@      �?             @        ������������������������       �                     �?        o       p                     @�q�q�?             @        ������������������������       �                     �?        q       r                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        t       �                   P`@��S�ۿ?8            �V@        u       �                    �?�*/�8V�?            �G@       v       {                    �?�>4և��?             <@        w       x                    �J@և���X�?             @        ������������������������       �                      @        y       z                   @_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        |                          j@�����?             5@        }       ~                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�X�<ݺ?             2@        �       �                   Xq@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �                     3@        �       �       
             �? qP��B�?            �E@       �       �                    �?г�wY;�?             A@        ������������������������       �                     $@        �       �                   Pa@ �q�q�?             8@        ������������������������       �                     "@        �       �                   �p@��S�ۿ?             .@       ������������������������       �                      @        �       �                   `b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?�"w����?2             S@       ������������������������       �        *             P@        �       �                    �?�8��8��?             (@        ������������������������       �                      @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��"�ű�?�            �i@        �       �                    �?�Pf����?9            �W@        �       �                   0d@�C��2(�?             6@       �       �                 @33�?8�Z$���?
             *@       �       �       
             �?      �?              @       �       �                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �c@�;�vv��?*            @R@        �       �                   �Z@���N8�?	             5@        ������������������������       �                      @        �       �                    S@�S����?             3@       �       �                    �?     ��?             0@       �       �                    �L@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�E��
��?!             J@       �       �                   `\@�θ�?            �C@        �       �                 @33�?      �?              @       �       �                   p`@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @`Jj��?             ?@       ������������������������       �                     =@        ������������������������       �                      @        �       �                   �p@$�q-�?             *@        �       �                   �n@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?�2����?M            �[@       �       �                   @E@���!pc�?'            �K@        �       �                   @^@ףp=
�?             $@        �       �                   `]@      �?             @        ������������������������       �                      @        �       �                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @a@�r����?            �F@       �       �                    �?@4և���?             <@       ������������������������       �                     7@        �       �                   0c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �N@������?             1@       �       �                    �?�	j*D�?             *@       �       �                    �L@�q�q�?
             (@       �       �                    @H@���!pc�?	             &@       �       �                    �F@���Q��?             @       �       �                    �D@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 pff�?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pt@�1�`jg�?&            �K@       �       �                   @[@�O4R���?%            �J@        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        "             I@        ������������������������       �                      @        �       �                 `ff�?`	�<��?^            �a@       �       �                    �?P�R�`M�?W            ``@        �       �                    �L@�eP*L��?             6@       �       �                    @H@�t����?	             1@        �       �                   �\@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �g@����q�?J            @[@       ������������������������       �        I            �Z@        ������������������������       �                      @        �       �                   d@�z�G��?             $@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�   Np	�?���Gw{�?<4WV���?�e��#��?5l7˓��?�$2���?UUUUUU�?UUUUUU�??4և���?�r
^N��?۶m۶m�?�$I�$I�?      �?      �?              �?      �?        333333�?ffffff�?�q�q�?9��8���?�������?333333�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�Q����?��Q���?B{	�%��?/�����?              �?y�5���?Cy�5��?UUUUUU�?UUUUUU�?r�q��?�q�q�?      �?      �?              �?      �?        �������?333333�?              �?      �?                      �?              �?d!Y�B�?ӛ���7�?�������?333333�?      �?                      �?              �?!Y�B�?��Moz��?9��8���?�q�q�?�������?�������?      �?      �?      �?                      �?              �?]t�E�?F]t�E�?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?                      �?y�5���?Cy�5��?;�;��?vb'vb'�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?XG��).�?��:��?b�a��?�y��y��?              �?�$I�$I�?۶m۶m�?vb'vb'�?�N��N��?      �?        Y�B��?zӛ����?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?              �?              �?Ũ�oS��?���u��?              �?�}�K�`�?C��6�S�?      �?      �?              �?d!Y�B�?Nozӛ��?�?xxxxxx�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�?�������?m�w6�;�?r1����?�m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?�a�a�?=��<���?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?��8��8�?      �?      �?              �?      �?                      �?              �?�}A_З?��}A�?�?�?              �?UUUUUU�?�������?              �?�?�������?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?(�����?Cy�5��?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ��q9�?�Ѹ���?�-q����?a�+F�?]t�E�?F]t�E�?;�;��?;�;��?      �?      �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ����Ǐ�?�8�?��y��y�?�a�a�?      �?        ^Cy�5�?(������?      �?      �?t�E]t�?F]t�E�?              �?      �?                      �?              �?;�;��?��؉���?ى�؉��?�؉�؉�?      �?      �?UUUUUU�?�������?      �?                      �?              �?���{��?�B!��?      �?                      �?;�;��?�؉�؉�?�������?�������?              �?      �?                      �?��7�}��?� O	��?F]t�E�?t�E]t�?�������?�������?      �?      �?              �?      �?      �?              �?      �?                      �?�������?�?n۶m۶�?�$I�$I�?      �?        333333�?�������?      �?                      �?xxxxxx�?�?vb'vb'�?;�;��?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?333333�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?�������?UUUUUU�?      �?                      �?              �?      �?              �?        A��)A�?�־a�?:�&oe�?�x+�R�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?o����?E�)͋?�?�	)y��?ձ�6Ls�?t�E]t�?]t�E�?�������?�������?�$I�$I�?�m۶m��?              �?      �?              �?                      �?���%�i�?�,�M�ɒ?      �?                      �?333333�?ffffff�?�q�q�?9��8���?              �?�������?333333�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��B�;         j                    �?6������?�           ��@               =                    �?J����*�?�            @v@                                  `@�����H�?�            `n@                                   �?���|���?             F@                                 `T@�חF�P�?             ?@                                   ^@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        	       
                    �? ��WV�?             :@       ������������������������       �                     3@                                  �^@؇���X�?             @       ������������������������       �                     @                                `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?8�Z$���?             *@        ������������������������       �                     �?                                   �?�8��8��?             (@                     
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  `Q@������?�            �h@                                  �a@      �?              @        ������������������������       �                     @                                   �J@�q�q�?             @        ������������������������       �                     �?                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               :                 ���@8��$��?|            �g@               %                    �?�	�(�Z�?z            �g@        !       "                   �d@z�G�z�?             $@       ������������������������       �                     @        #       $                     J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        &       -                    @L@@]����?u            @f@       '       ,                   @[@@�`%���?`            `b@        (       +                    c@�����H�?             "@        )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        Z            @a@        .       1                   �i@��� ��?             ?@        /       0                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        2       7                   ht@HP�s��?             9@       3       6                    �L@���N8�?             5@        4       5                   Hp@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        8       9                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ;       <                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        >       E                   `d@�������?B            @\@        ?       D                   �e@��� ��?             ?@       @       C                    �? 	��p�?             =@        A       B                    `Q@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                      @        F       O                    �?v�2t5�?1            �T@        G       H                    �?��2(&�?             6@        ������������������������       �                     &@        I       N       	             �?���!pc�?             &@        J       M                    @K@���Q��?             @       K       L                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        P       i                   (u@      �?$             N@       Q       h                   �n@���y4F�?#            �L@       R       g       	             �?և���X�?             <@       S       T                 ����?�q�q�?             8@        ������������������������       �                     @        U       Z                   b@��.k���?             1@        V       W                 ����?z�G�z�?             @        ������������������������       �                     @        X       Y                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        [       `                   �k@�q�q�?             (@        \       _                    �?���Q��?             @       ]       ^                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        a       f                    �?؇���X�?             @       b       c                   �l@r�q��?             @        ������������������������       �                     @        d       e                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        ������������������������       �                     @        k       �                    �?d}h���?�            �w@        l       �                    �?6�\"���?R            �_@       m       �                 ����?�'�=z��??            �X@        n                           �?�3Ea�$�?             G@       o       p                   �`@(L���?            �E@       ������������������������       �                     8@        q       |                    �?�����?             3@       r       {                    m@      �?	             0@       s       z                   �b@�q�q�?             (@       t       y                   �b@z�G�z�?             $@       u       v                    @K@�q�q�?             @        ������������������������       �                     @        w       x                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        }       ~                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �F@Ȩ�I��?#            �J@        ������������������������       �                      @        �       �                    �?f.i��n�?            �F@        �       �                    �?j���� �?             1@       �       �                   �Z@���!pc�?             &@        ������������������������       �                      @        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                    `P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                   `_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @؇���X�?             <@       �       �                   �t@�<ݚ�?             2@       �       �                 `ff�?@�0�!��?             1@       �       �                    c@@4և���?
             ,@       ������������������������       �                     &@        �       �                   `^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?      �?             <@        ������������������������       �                     @        �       �                 `ff @�q�q�?             5@       �       �                   @f@�d�����?             3@       �       �                    �?@�0�!��?             1@        �       �                   xq@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �[@@4և���?	             ,@        �       �                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��<VO�?�            `o@       �       �                    �?�c:��?w             g@       �       �                    b@���Hx�?[             b@        ������������������������       �                     7@        �       �                    @Q@����W1�?K            @^@       �       �                    �?2Tv���?J             ^@       �       �                    �?Ĝ�oV4�?9            �V@        �       �                 ����?������?             1@       �       �                   `c@      �?              @       �       �                   �a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�����?.            �R@        �       �                 ����?@4և���?             <@       ������������������������       �        
             2@        �       �                     G@z�G�z�?             $@        �       �                    ]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @�q��/��?             G@       �       �                   0c@��hJ,�?             A@       �       �                    �O@     ��?             @@       �       �                   �\@`Jj��?             ?@        �       �                   @a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �Z@ 	��p�?             =@        �       �                 033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     :@        ������������������������       �                     �?        ������������������������       �                     D@        �       �                    �J@��v����?'            �P@        �       �                   Pm@�	j*D�?	             *@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@       �       �                    Z@      �?              @        ������������������������       �                     @        �       �                    @z�G�z�?             @       �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �_@h�WH��?             K@       �       �                 ����?�?�|�?            �B@        �       �                   �]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @@        �       �                    �O@������?
             1@       ������������������������       �                     $@        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��X�5�?��S�$e�?mjS����?%+Y�JV�?�q�q�?�q�q�?]t�E]�?F]t�E�?�Zk����?��RJ)��?�������?�������?      �?                      �?O��N���?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?              �?�n-;�?���/M�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?vX�Q�}�?�x��* �?������?L� &W�?�������?�������?      �?              �?      �?              �?      �?        �g<��?�as�Ü?���E��?���+�{?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?        �{����?�B!��?UUUUUU�?UUUUUU�?              �?      �?        q=
ףp�?{�G�z�?��y��y�?�a�a�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�ZX驅�?��S+=�?�B!��?�{����?�{a���?������?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?        �ڕ�]��?��+Q��?��.���?t�E]t�?      �?        F]t�E�?t�E]t�?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?(������?6��P^C�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?�?�������?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?      �?                      �?      �?        ۶m۶m�?I�$I�$�?O���t:�?Y,��b�?|��|�?|���?����7��?��,d!�?⎸#��?w�qG��?      �?        Q^Cy��?^Cy�5�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�	�[���?+�R��?              �?�>�>��?�`�`�?�������?ZZZZZZ�?F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?۶m۶m�?�q�q�?9��8���?�������?ZZZZZZ�?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?y�5���?Cy�5��?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        �ZEtJu�?�Tw�V�?8��Moz�?Y�B���?9��8��?9��8���?              �?���|���?��eP*L�?�������?�������?����?�!�!�?�?xxxxxx�?      �?      �?�������?�������?      �?                      �?              �?              �?v�)�Y7�?�Ϻ���?�$I�$I�?n۶m۶�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?��Mozӻ?�B����?�������?KKKKKK�?      �?      �?�B!��?���{��?�������?333333�?      �?                      �?              �?      �?              �?                      �?�{a���?������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?*g��1�?5&����?;�;��?vb'vb'�?              �?�q�q�?r�q��?      �?      �?              �?�������?�������?      �?      �?      �?                      �?      �?                      �?B{	�%��?��^B{	�?к����?*�Y7�"�?�������?�������?              �?      �?                      �?�?xxxxxx�?              �?�$I�$I�?۶m۶m�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�7         H                   P`@U�ք�?�           ��@               3                   P`@j=M>�:�?�            �s@               .       	             �?��+7��?X            @a@              %                    �?HC>���?P            �^@                                 `_@p���p�?@            �Y@                                 `[@�����?(            �P@        ������������������������       �                     6@                                   �?��S�ۿ?            �F@        	       
                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @                      
             �?��Y��]�?            �D@                                 `_@P�Lt�<�?             C@       ������������������������       �                     >@                                   �K@      �?              @       ������������������������       �                     @                                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �]@tk~X��?             B@                                  �?HP�s��?             9@                                  `@ �q�q�?             8@                                   @M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?                                    �?�eP*L��?             &@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        !       "                    �L@����X�?             @        ������������������������       �                     @        #       $                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        &       )                    �?�����?             3@       '       (                   (r@�C��2(�?	             &@       ������������������������       �                     $@        ������������������������       �                     �?        *       -                    �?      �?              @       +       ,                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        /       0                    �?     ��?             0@        ������������������������       �                     "@        1       2                    `@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        4       ?                    �?��/eA��?h             f@        5       8                 033�?��c:�?             G@       6       7                    �?���N8�?             5@        ������������������������       �                     @        ������������������������       �                     0@        9       >                 `ff@H%u��?             9@       :       ;       	             �?�nkK�?             7@       ������������������������       �        	             1@        <       =                    �K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        @       A                   0q@�z�N��?M            ``@       ������������������������       �        <             Y@        B       G                    �?��a�n`�?             ?@       C       D                    �?XB���?             =@       ������������������������       �                     ;@        E       F                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        I       �                    �?@<QR���?           0z@       J       �                    �?��<b���?�            �o@       K       R                    I@b<g���?�            `k@        L       Q                    �?      �?              @       M       N                    \@����X�?             @        ������������������������       �                     �?        O       P                    `@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        S       �                    �P@�$
��
�?�            `j@       T       }                   h@<��u���?�            `i@       U       b                    �?P���+�?�            �h@       V       W                   pl@x�C����?d            �b@        ������������������������       �        1            �Q@        X       Y                    �?XI�~�?3            @S@        ������������������������       �                     <@        Z       [                    @G@ i���t�?"            �H@       ������������������������       �                     :@        \       ]                   �\@��<b���?             7@        ������������������������       �                     @        ^       _                    @L@�}�+r��?             3@       ������������������������       �        	             (@        `       a                 @33�?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        c       r       	             �?ҳ�wY;�?            �I@       d       i                 ����?�eP*L��?            �@@       e       f                   `j@����X�?
             ,@        ������������������������       �                     @        g       h                     O@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        j       q                    `@�d�����?	             3@       k       l                   �k@�eP*L��?             &@        ������������������������       �                     @        m       n                     H@      �?              @        ������������������������       �                     @        o       p                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        s       |                   d@r�q��?
             2@       t       {                    �?      �?             (@       u       v                   �\@"pc�
�?             &@        ������������������������       �                     �?        w       x                    �?ףp=
�?             $@        ������������������������       �                     @        y       z                   pn@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ~                          pn@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�ʻ����?             A@       �       �                    �?     ��?             @@        �       �                    p@      �?	             0@       �       �                    @J@�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                    �M@z�G�z�?             @        ������������������������       �                      @        �       �                 lffֿ�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �O@     ��?	             0@       �       �                    �?d}h���?             ,@       ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�)��V��?m            �d@       �       �                    s@���Q��?:            �W@       �       �                 ����?k��9�?7            �V@       �       �                    P@�ɞ`s�?&            �N@        ������������������������       �                     @        �       �                    �?�d�����?#            �L@       �       �                   0d@�#-���?            �A@       ������������������������       �                     :@        �       �                    �?�q�q�?             "@       �       �                    a@      �?              @       ������������������������       �                     @        �       �                    �?      �?             @       �       �                   l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `\@�eP*L��?             6@        �       �                    m@      �?              @       ������������������������       �                     @        �       �                   �[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?և���X�?             ,@       �       �                    �?���|���?             &@        �       �                   d@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �J@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   `e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �U@J�8���?             =@        ������������������������       �                     @        �       �                   �d@R�}e�.�?             :@        �       �                    �?�q�q�?             "@       �       �                 033�?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�IєX�?
             1@        ������������������������       �                      @        �       �                   Pm@�����H�?             "@       ������������������������       �                     @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?��UV�?3            �Q@        �       �                    �?���7�?             6@       ������������������������       �                     4@        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ZՏ�m|�?%            �H@        �       �                   �a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �m@��p\�?            �D@       �       �                    �?�����H�?             ;@       �       �                   �`@d}h���?             ,@       �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                   �h@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     ,@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ᓔ��?�5�;��?y�y��?�����?Y�B��?zӛ����?�y��!�?�!XG���?C��ڸ?�E|���?���@��?g��1��?              �?�?�������?      �?      �?      �?                      �?������?8��18�?(�����?���k(�?              �?      �?      �?              �?      �?      �?      �?                      �?              �?9��8���?r�q��?{�G�z�?q=
ףp�?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        ]t�E�?t�E]t�?      �?      �?              �?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?Q^Cy��?^Cy�5�?]t�E�?F]t�E�?      �?                      �?      �?      �?333333�?�������?      �?                      �?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        Cr��ѿ?��
��?�7��Mo�?-d!Y��?�a�a�?��y��y�?              �?      �?        ���Q��?)\���(�?d!Y�B�?�Mozӛ�?              �?UUUUUU�?�������?      �?                      �?      �?        ձ�6Ls�?qBJ�eD�?              �?�c�1Ƹ?�s�9��?�{a���?GX�i���?              �?      �?      �?              �?      �?              �?        �8�)�?\��+��?��,d!�?��Moz��?֫W�^��?�P�B�
�?      �?      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?              �?        =:�oL�??�A��?��P@���?�)���d�?���/M�?�Q7���?�n0E>��?���L�?      �?        5�wL��?V~B����?      �?        /�����?����X�?      �?        ��,d!�?��Moz��?              �?�5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?      �?                      �?�������?�������?t�E]t�?]t�E�?�$I�$I�?�m۶m��?      �?        F]t�E�?]t�E�?              �?      �?        Cy�5��?y�5���?t�E]t�?]t�E�?              �?      �?      �?      �?              �?      �?              �?      �?              �?        �������?UUUUUU�?      �?      �?/�袋.�?F]t�E�?              �?�������?�������?      �?        ۶m۶m�?�$I�$I�?      �?                      �?              �?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?<<<<<<�?�������?      �?      �?      �?      �?9��8���?�q�q�?              �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?              �?      �?۶m۶m�?I�$I�$�?              �?      �?              �?              �?        GS��r�?]V��F�?333333�?�������?�'}�'}�?[�[��?mާ�d�?&C��6��?              �?Cy�5��?y�5���?�A�A�?_�_�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?      �?              �?      �?                      �?      �?        ]t�E�?t�E]t�?      �?      �?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?]t�E]�?F]t�E�?333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        |a���?�rO#,��?      �?        �;�;�?'vb'vb�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?�?�?              �?�q�q�?�q�q�?              �?      �?      �?              �?      �?              �?        6��9�?2~�ԓ��?F]t�E�?�.�袋�?              �?      �?      �?      �?                      �?9/����?�>4և��?      �?      �?      �?                      �?��+Q��?�]�ڕ��?�q�q�?�q�q�?۶m۶m�?I�$I�$�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��B�;         �                    �?0����?�           ��@              %                    �?��YB�8�?           �y@                                   �J@TV����?*            �M@                                   �?����X�?             5@                                 xq@���y4F�?             3@                                 �Q@      �?             0@        ������������������������       �                     �?                      
             �?��S�ۿ?             .@        	                            H@z�G�z�?             @        
                           `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                   �?�q�q�?             @        ������������������������       �                     �?                                  �s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �?p9W��S�?             C@                                   �?      �?
             (@                                 �Z@"pc�
�?	             &@                      
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?               $                    �?$�q-�?             :@                                  �?      �?	             0@        ������������������������       �                      @                #                   �s@      �?              @       !       "                   `^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        &       u                    �?��g�g�?�             v@       '       l                   Ps@ȵHPS!�?�            �q@       (       9                    @G@8�����?�            �p@        )       4       	             �?Jm_!'1�?            �H@       *       1       
             �?������?            �D@       +       ,                   �m@�}�+r��?             C@       ������������������������       �                     6@        -       0                    �?      �?	             0@        .       /                   pb@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        2       3                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        5       6                    �B@      �?              @        ������������������������       �                      @        7       8                     @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        :       E                   i@<�*/�{�?�             k@        ;       @       
             �?��F�D�?9            �X@       <       =                    �? �)���?.            @T@       ������������������������       �                    �M@        >       ?                   �_@���7�?             6@        ������������������������       �                     �?        ������������������������       �                     5@        A       B                    �N@�X�<ݺ?             2@       ������������������������       �                     *@        C       D                   `a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        F       G                   @i@�^����?K            �]@        ������������������������       �                     �?        H       c       
             �?�����H�?J            @]@       I       ^       	             �?W�!?�?=            �X@       J       ]                   �b@|)����?7            �V@       K       \                    �?���M�?5            @V@       L       U                    �?���}<S�?(            @Q@        M       N                    �?"pc�
�?             6@        ������������������������       �                      @        O       P                   �i@ףp=
�?             4@        ������������������������       �                     �?        Q       T                   �`@�}�+r��?
             3@        R       S                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        V       [                   �[@`�q�0ܴ?            �G@        W       X                   �Z@�����H�?	             2@       ������������������������       �                     ,@        Y       Z                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     4@        ������������������������       �                      @        _       b                    �?      �?              @        `       a                   �d@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        d       e                   �l@r�q��?             2@       ������������������������       �                     $@        f       i                 033�?      �?              @        g       h                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        j       k                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        m       n                    �?���Q��?             4@        ������������������������       �                     @        o       t                    �?z�G�z�?
             .@       p       q                    T@      �?             (@        ������������������������       �                      @        r       s                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        v       �                    �?@�0�!��?,             Q@        w       x                    �K@�n_Y�K�?             :@        ������������������������       �                     @        y       �                    �O@z�G�z�?             4@       z       {       
             �?$�q-�?	             *@        ������������������������       �                     @        |                        ����?r�q��?             @        }       ~                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     P@և���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���N8�?             E@        ������������������������       �                     @        �       �                   �Z@�X�<ݺ?             B@        ������������������������       �                      @        ������������������������       �                     A@        �       �                   @E@�f,0Bo�?�            t@        �       �                    �L@p�ݯ��?             C@       �       �                   �?���y4F�?             3@        �       �                    �?X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�\��N��?             3@       �       �       	             �?�q�q�?	             .@       �       �                    �M@�q�q�?             (@        ������������������������       �                     @        �       �                    �?      �?              @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?l�?����?�            �q@       �       �                    @pŰ�e��?�            �h@       �       �                    �?��~F�<�?�            �h@       �       �                    �?�s0jo�?z            `g@        ������������������������       �        !             G@        �       �                    �?�lm�9�?Y            �a@        ������������������������       �                    �D@        �       �       	             �?`2U0*��?@             Y@        �       �                 ����?��(\���?             D@       �       �                   �s@��a�n`�?             ?@       �       �                   @[@��S�ۿ?             >@        ������������������������       �                      @        ������������������������       �                     <@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �_@ �.�?Ƞ?'             N@        �       �                   �o@ ��WV�?             :@       ������������������������       �                     4@        �       �                   `p@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     A@        �       �                    p@z�G�z�?             $@       �       �                   0`@      �?              @        ������������������������       �                     @        �       �                   �h@�q�q�?             @        ������������������������       �                     �?        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    _@����X�?3             U@        �       �                   �q@"pc�
�?            �@@       �       �                    �?ףp=
�?             >@       �       �                   �c@      �?             8@       �       �                    �?      �?             (@       �       �                   �o@ףp=
�?             $@       ������������������������       �                     @        �       �                   �p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     @        �       �                    s@ҳ�wY;�?            �I@       �       �                    �?�K��&�?            �E@        �       �                   �c@      �?             6@       �       �                 ����?b�2�tk�?             2@       �       �                   �_@���|���?             &@        ������������������������       �                     @        �       �                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����?�q�q�?             5@       �       �                    `@8�Z$���?
             *@        ������������������������       �                     �?        �       �                   pf@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                 ����?      �?              @        ������������������������       �                     �?        �       �                    b@և���X�?             @       �       �                   �k@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B�  ���^L�?���Y�?��]=�?V�����?u_[4�?E�pR���?�m۶m��?�$I�$I�?6��P^C�?(������?      �?      �?              �?�������?�?�������?�������?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?l(�����?�k(����?      �?      �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?;�;��?�؉�؉�?      �?      �?              �?      �?      �?      �?      �?      �?                      �?              �?              �?��}ylE�?ي����?�؉�؉�?��N��N�?���f�?�τ?��?������?����X�?������?�|����?(�����?�5��P�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�������?UUUUUU�?      �?                      �?��K�%�?��G���?[�R�֯�?j�J�Z�?�����H�?X�<ݚ�?              �?F]t�E�?�.�袋�?      �?                      �?�q�q�?��8��8�?              �?�������?�������?              �?      �?        W'u_�?u_[4�?      �?        �q�q�?�q�q�?1ogH�۹?�v���?h�h��?��/��/�?�E(B�?��^����?d!Y�B�?ӛ���7�?F]t�E�?/�袋.�?      �?        �������?�������?      �?        (�����?�5��P�?      �?      �?      �?                      �?              �?W�+�ɥ?��F}g��?�q�q�?�q�q�?              �?      �?      �?      �?                      �?              �?              �?      �?              �?      �?�������?333333�?      �?                      �?              �?UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?�������?333333�?      �?        �������?�������?      �?      �?      �?        �������?�������?      �?                      �?              �?�������?ZZZZZZ�?ى�؉��?;�;��?      �?        �������?�������?;�;��?�؉�؉�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?              �?      �?                      �?�a�a�?��y��y�?              �?�q�q�?��8��8�?      �?                      �?����j�?���+�T�?Cy�5��?^Cy�5�?(������?6��P^C�?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?      �?                      �?              �?y�5���?�5��P�?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?hw4�a�?ƿD\n�?���a���?gв�9��?�;�Y�?&���0�?Q9"�P�?�и[�?      �?        ���S��?t�n���?      �?        ���Q��?{�G�z�?�������?333333�?�s�9��?�c�1Ƹ?�������?�?              �?      �?                      �?      �?        wwwwww�?�?O��N���?;�;��?      �?        �������?UUUUUU�?              �?      �?              �?        �������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?              �?�m۶m��?�$I�$I�?/�袋.�?F]t�E�?�������?�������?      �?      �?      �?      �?�������?�������?      �?              �?      �?              �?      �?                      �?      �?              �?                      �?�������?�������?��)kʚ�?���)k��?      �?      �?9��8���?�8��8��?]t�E]�?F]t�E�?              �?      �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKǅ�h��B�1         V                    �?�+	G�?�           ��@               ;                    �?~)6ź��?�            �u@                                 @E@Ĝ�oV4�?�            q@                      	             �?�q�q�?             8@              
                   @^@      �?             4@                                ����?X�<ݚ�?             "@        ������������������������       �                     @               	                   �]@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @               :                   �g@0*��ɾ?�             o@              -                   �a@Pi�M`�?�            �n@              ,                 ���@�m��1�?�             j@              +                   Pd@�:���ΰ?~            �i@                                  @L@��vp(�?W            �a@                                 �[@���͡?C            @\@                                   @H@؇���X�?	             ,@                                  �?      �?              @                     
             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        :            �X@               *                    �?�>4և��?             <@              )       
             �?��<b���?             7@                                @33�?      �?             4@        ������������������������       �                      @        !       (                    �?�q�q�?             (@       "       %                 ����?�eP*L��?             &@       #       $                   @`@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        &       '                    �P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        '            @P@        ������������������������       �                      @        .       9                   �f@�ݜ�?            �C@       /       4                   �b@�KM�]�?             C@        0       1                   `_@�q�q�?             "@        ������������������������       �                      @        2       3                   �m@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        5       6                   �r@XB���?             =@       ������������������������       �                     :@        7       8                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        <       U                    �?؀�:M�?-            �R@       =       B                    �?��T���?,            @R@        >       A                   �a@�r����?             .@        ?       @       	             �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        C       F                    �?>���Rp�?%             M@       D       E                    �R@(;L]n�?             >@       ������������������������       �                     =@        ������������������������       �                     �?        G       T                   `c@���>4��?             <@       H       S                   pk@�ՙ/�?             5@       I       R                    �O@��S���?	             .@       J       K                     M@���|���?             &@        ������������������������       �                      @        L       Q                    �?�<ݚ�?             "@       M       N                    �M@      �?              @        ������������������������       �                      @        O       P                   �V@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        W       �       	             �?f�g��N�?�            0x@       X       �                    �?<+̫���?�            Pv@        Y       |                    �?l�Ӑ���?9            �U@       Z       e                    �?p�EG/��?'            �O@        [       \                   `X@�d�����?             3@        ������������������������       �                     @        ]       d                    c@      �?
             0@       ^       _       
             �?��S�ۿ?	             .@        ������������������������       �                      @        `       a                   0e@$�q-�?             *@       ������������������������       �                      @        b       c                   �l@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        f       o                    �?      �?             F@       g       h                   0b@H%u��?             9@       ������������������������       �        
             1@        i       j                 `ff�?      �?              @        ������������������������       �                     @        k       l                   Pb@���Q��?             @        ������������������������       �                      @        m       n                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        p       q                    �L@D�n�3�?             3@        ������������������������       �                     @        r       y                    �?������?             .@       s       x                 ����?"pc�
�?             &@        t       u                    `P@�q�q�?             @        ������������������������       �                     �?        v       w                   c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        z       {                   c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        }       �                    �?      �?             8@       ~                           @F@z�G�z�?             .@        ������������������������       �                     �?        �       �                    \@؇���X�?             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?             *@        ������������������������       �                     @        �       �                     N@      �?              @        �       �                   �l@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �Q@���?�            �p@       �       �                    �?�ƫ�%�?�            �p@       �       �                   �e@�n����?�            �i@       �       �                    c@��Y��]�?�            �i@       �       �                 ����? S5W�?v             g@        �       �                   P`@`���i��?             F@       ������������������������       �                     ?@        �       �                   �`@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        Z            �a@        �       �                    �?z�G�z�?             4@       �       �                   �j@"pc�
�?             &@        ������������������������       �                     @        �       �                   �n@����X�?             @        ������������������������       �                     �?        �       �                   xu@r�q��?             @       ������������������������       �                     @        �       �                   pc@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        �       �                    �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ����?�r����?%             N@        �       �                    �?R�}e�.�?             :@        �       �                   �`@      �?             ,@       �       �                    �?�z�G��?             $@        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                   `\@г�wY;�?             A@        �       �                    �L@؇���X�?             @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?��S���?             >@       �       �                    �?������?             1@        ������������������������       �                     @        �       �                    �?���Q��?             $@        �       �                 433�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?$�q-�?             *@       ������������������������       �                     $@        �       �                    p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  ��C�l�?z?+^���?>��h���?��\&$�?�!�!�?����?�������?�������?      �?      �?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?�>���?��G
&s�?����/�?S���.�?ى�؉��?vb'vb'�?�~�����?�H%�e�?z�'Ni�?f��k�?$��Co�?x�!���?۶m۶m�?�$I�$I�?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?              �?        �$I�$I�?�m۶m��?��,d!�?��Moz��?      �?      �?      �?        �������?�������?t�E]t�?]t�E�?�m۶m��?�$I�$I�?              �?      �?              �?      �?              �?      �?              �?              �?              �?              �?                      �?\��[���?�i�i�?�k(���?(�����?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?              �?      �?        GX�i���?�{a���?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?v�)�Y7�?E>�S��?�z��ի�?�B�
*�?�������?�?333333�?�������?              �?      �?              �?        GX�i���?�i��F�?�?�������?              �?      �?        n۶m۶�?I�$I�$�?�<��<��?�a�a�?�������?�?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?      �?      �?        �������?UUUUUU�?              �?      �?                      �?              �?      �?                      �?      �?        �D�f�.�?��]&B4�? D�D��?|W|W�?/�I���?�7[�~��?Y�eY�e�?�4M�4M�?Cy�5��?y�5���?              �?      �?      �?�������?�?      �?        �؉�؉�?;�;��?      �?        �������?�������?      �?                      �?              �?      �?      �?���Q��?)\���(�?              �?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        (������?l(�����?      �?        �?wwwwww�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?      �?�������?�������?      �?        �$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?t��:W�?��oS��?�as�ì?��x�3�?j6��bP�?�<����?������?8��18�?@bw�#v?<����?F]t�E�?F]t�E�?              �?;�;��?�؉�؉�?      �?                      �?              �?�������?�������?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?9��8���?              �?      �?      �?              �?      �?              �?        �?�������?�;�;�?'vb'vb�?      �?      �?333333�?ffffff�?      �?              �?      �?      �?                      �?      �?                      �?�?�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�?xxxxxx�?�?      �?        333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         `                 ����?6������?�           ��@              -                    �?��v��?�            �w@              ,                   �g@Ί�C�o�?�            �o@                                 �Y@� ��?�             o@                      	             �?"pc�
�?             &@                                  �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        	       
                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �c@��w\ud�?�            �m@                                   �?D�n�3�?             3@        ������������������������       �                      @        ������������������������       �                     &@                                  �n@����1�?�            `k@                                  �?0Ƭ!sĮ?X             `@                      
             �?���y4F�?             3@        ������������������������       �                     $@                                  �d@X�<ݚ�?             "@                                 �m@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        M            �[@               '                    �?>���a��?5            �V@              $                    @O@Х-��ٹ?-            �R@                                  �?�\=lf�?(            �P@        ������������������������       �                     5@               #                   �b@��<b�ƥ?             G@               "       
             �?�IєX�?
             1@               !                   �a@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        %       &                 ����?      �?              @        ������������������������       �                     @        ������������������������       �                     @        (       )                    @O@�r����?             .@       ������������������������       �                     &@        *       +                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        .       _                   �f@-"� ��?U            ``@       /       @                   �i@PlX=��?R            �_@        0       ?                    @N@�z�6�?&             O@       1       2                    �?����|e�?              K@       ������������������������       �                     @@        3       <                    �?8�A�0��?             6@       4       ;                   �b@��S���?
             .@       5       :                   @E@���!pc�?             &@        6       9                    �?���Q��?             @       7       8                    �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        =       >                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        A       F                    �?��
ц��?,            @P@        B       E                    �?     ��?             0@       C       D                    �J@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        G       T                    �?Tt�ó��?!            �H@        H       S                    �?��}*_��?             ;@       I       P                   �b@��s����?             5@       J       K                    �?�����H�?
             2@       ������������������������       �                     (@        L       O                   �d@�q�q�?             @       M       N                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Q       R                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        U       ^                    �?�GN�z�?             6@       V       W                   �_@�q�q�?             .@        ������������������������       �                     @        X       [                   @l@X�<ݚ�?             "@        Y       Z                   `^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        \       ]                 ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        a       |                    a@x�����?�            �u@        b       c                   �]@��(\���?5             T@        ������������������������       �                     ;@        d       m                    ^@���C��?$            �J@        e       j                    �?      �?              @       f       i                 033�?z�G�z�?             @       g       h                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        k       l                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        n       u                    �?��S�ۿ?            �F@       o       p                 `ff�?г�wY;�?             A@       ������������������������       �                     3@        q       t                   �`@��S�ۿ?	             .@        r       s                   0`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        v       w                 ����?"pc�
�?             &@       ������������������������       �                     @        x       {                    @���Q��?             @       y       z                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        }       �                    �?��v4Ք�?�            �p@        ~       �                    �?      �?<            �V@              �                   �s@�v:���?,             Q@       �       �                   �`@�ɞ`s�?)            �N@       �       �                   �l@      �?             @@        �       �                    `P@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   p@����X�?             5@       �       �                    @      �?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                   @_@�C��2(�?             &@       ������������������������       �                      @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     K@ܷ��?��?             =@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   �o@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �? �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?؇���X�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?�C��2(�?             6@        �       �                   0i@"pc�
�?             &@        ������������������������       �                     @        �       �                   �_@�q�q�?             @       ������������������������       �                     @        �       �                 033�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 ����?l�oA�?x            �f@        �       �                   �k@�BbΊ�?$             M@        ������������������������       �                     &@        �       �                    �?(���@��?            �G@        �       �                    �M@�z�G��?             $@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���@��?            �B@        ������������������������       �                     @        �       �                 ����?r٣����?            �@@       �       �                    �?������?             >@       �       �                   pl@l��
I��?             ;@        ������������������������       �                     @        �       �                    �?��2(&�?             6@       ������������������������       �        	             ,@        �       �                   `]@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@������?T            �^@       �       �                   pa@t�e�í�?.            �P@       �       �                   `_@�X�<ݺ?%             K@        �       �                     P@�8��8��?             8@       �       �                   po@�nkK�?             7@       ������������������������       �        
             ,@        �       �                   �_@�����H�?             "@       �       �                   pp@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �J@(;L]n�?             >@        �       �                   @_@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?8�Z$���?	             *@       �       �                   �p@z�G�z�?             $@       ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �R@�h����?&             L@       ������������������������       �        %            �K@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  ��X�5�?��S�$e�?&���P��?���>^�?�,˲,��?5M�4M��?q����?<v5,���?F]t�E�?/�袋.�?�q�q�?�q�q�?              �?      �?              �?      �?              �?      �?        �����?�z1�z1�?l(�����?(������?              �?      �?        �Ν;w��?Ĉ#F��?����?����?6��P^C�?(������?      �?        r�q��?�q�q�?�������?�������?              �?      �?              �?              �?        J��I���?؂-؂-�?K~��K�?O贁N�?"=P9���?g��1��?      �?        ��7��M�?d!Y�B�?�?�?]t�E�?F]t�E�?      �?                      �?      �?              �?              �?      �?              �?      �?        �?�������?              �?      �?      �?      �?                      �?              �?�U���g�?ձ�6L�?��`0�?�|>����?�Zk����?J)��RJ�?	�%����?����K�?              �?颋.���?/�袋.�?�?�������?F]t�E�?t�E]t�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?              �?�;�;�?�؉�؉�?      �?      �?      �?      �?      �?                      �?      �?        /�����?h�����?_B{	�%�?B{	�%��?z��y���?�a�a�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?              �?]t�E�?�袋.��?UUUUUU�?UUUUUU�?              �?r�q��?�q�q�?      �?      �?              �?      �?        �������?�������?              �?      �?                      �?      �?        �A�A�?��o��o�?333333�?�������?              �?"5�x+��?\�琚`�?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�������?�?�?              �?�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?/�袋.�?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?G��f,�?.A�~�4�?      �?      �?�������?<<<<<<�?&C��6��?mާ�d�?      �?      �?]t�E�?F]t�E�?      �?                      �?�$I�$I�?�m۶m��?      �?      �?      �?                      �?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?a���{�?��=���?�������?333333�?              �?      �?      �?      �?                      �?UUUUUU�?�������?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        ]t�E�?F]t�E�?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ]��ҟ��?4O��I�?���=��?�{a��?              �?R�٨�l�?W�+���?ffffff�?333333�?      �?              �?      �?      �?                      �?к����?L�Ϻ��?              �?|���?>���>�?�?wwwwww�?h/�����?Lh/����?      �?        t�E]t�?��.���?              �?      �?      �?              �?      �?                      �?              �?������?p>�cp�?�rv��?�1����?�q�q�?��8��8�?UUUUUU�?UUUUUU�?d!Y�B�?�Mozӛ�?              �?�q�q�?�q�q�?�������?�������?      �?                      �?              �?      �?        �?�������?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?;�;��?;�;��?�������?�������?              �?�������?333333�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK텔h��B@;         v                    �?�Z���?�           ��@              O                    �?225,���?�            �v@                                 @E@�2�MA��?�            �q@               	                    �?�4�����?             ?@                                ����?�n_Y�K�?             *@                                 �b@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        
                        ����?�����H�?             2@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             (@               N                   h@     ��?�             p@              -                    @L@������?�            �o@              (                   �f@f�1�?z             g@                                  �?���fG��?t             f@                     	             �?@�z�G�?f             d@                                   �?������?/             R@                                 @[@h�����?$             L@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �j@@3����?"             K@                                ����?���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                     0@        ������������������������       �        7             V@                '       
             �?�t����?             1@        !       "                   �h@      �?              @        ������������������������       �                     �?        #       &                    @F@؇���X�?             @        $       %                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        )       ,                    �?      �?              @       *       +                    @C@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        .       G       
             �?���L��?(            �Q@       /       @                   `q@�	j*D�?             J@       0       1                    �L@      �?             D@        ������������������������       �                     @        2       =                    �?<ݚ)�?             B@       3       <                   Pd@J�8���?             =@       4       7                    �?�\��N��?             3@        5       6                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        8       ;                   �b@     ��?
             0@       9       :                   @n@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        >       ?                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        A       F                 @33�?�8��8��?             (@        B       C                    �?      �?              @        ������������������������       �                     @        D       E                   d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        H       I                    �?�X�<ݺ?             2@       ������������������������       �                     $@        J       K                   �k@      �?              @        ������������������������       �                     @        L       M                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        P       S                    �?      �?8             T@        Q       R                    �?      �?             0@       ������������������������       �                     ,@        ������������������������       �                      @        T       m                    �?      �?1             P@       U       l                   pq@����e��?            �@@       V       _                    �?���>4��?             <@        W       X                   `_@�<ݚ�?             "@        ������������������������       �                     @        Y       Z                    �?���Q��?             @        ������������������������       �                     �?        [       \                    �?      �?             @        ������������������������       �                     �?        ]       ^                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        `       k       	             �?D�n�3�?             3@       a       b                   �\@��S���?             .@        ������������������������       �                      @        c       j                 033�?�n_Y�K�?             *@       d       e                   �g@�eP*L��?	             &@        ������������������������       �                     @        f       g                   �o@����X�?             @        ������������������������       �                     @        h       i                   b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        n       u                   �r@��a�n`�?             ?@       o       t                     K@��S�ۿ?             >@        p       q                   �`@z�G�z�?             $@       ������������������������       �                     @        r       s                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        w       �                    �?p�5� ��?�            �v@        x       �                    �P@`��_��?+            �Q@       y       �       	             �?�eP*L��?(            �P@       z       �       
             �?      �?"             L@       {       �                   �`@v�X��?             F@        |                           �?      �?	             0@        }       ~                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@�	j*D�?             *@       �       �                    `@"pc�
�?             &@       �       �                   �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   pl@ �Cc}�?             <@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �k@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�}�+r��?             3@        �       �                   �x@z�G�z�?             @        ������������������������       �                      @        �       �                   pc@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             ,@        �       �                   �q@�q�q�?             (@       �       �                 ����?z�G�z�?             $@        ������������������������       �                     @        �       �                     H@      �?             @        ������������������������       �                     �?        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    d@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ȁZ|� �?�            �r@       �       �                   pa@��w"�"�?�            �n@       �       �                   �h@ ��^og�?u            �f@        ������������������������       �        5             U@        �       �                    �M@�"P��?@            �X@       �       �                    @M@ ����?,            @P@       �       �       	             �?�����?*            �O@       �       �                   �\@�8��8��?(             N@        �       �                    �?8�Z$���?             :@       �       �                   �Z@�}�+r��?             3@       ������������������������       �                     &@        �       �                    @K@      �?              @       ������������������������       �                     @        �       �                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                    @J@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �_@г�wY;�?             A@       �       �                   Pi@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     .@        �       �                   �n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   p`@г�wY;�?             A@        �       �                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@        �       �                   b@��f/w�?)            �N@        �       �                    �?�ՙ/�?             5@       �       �                   �_@�n_Y�K�?             *@       �       �                    �?؇���X�?             @       �       �                    �C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �d@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             D@        ������������������������       �                     1@        �       �                 ����?��<b���?             7@        ������������������������       �                     �?        �       �                     O@"pc�
�?             6@       �       �                    �?ףp=
�?             4@       ������������������������       �                     (@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �Z@���B���?"             J@        ������������������������       �                     @        �       �                    �?�*/�8V�?             �G@        �       �                    @G@�t����?             1@        ������������������������       �                      @        �       �                    �?z�G�z�?             .@       �       �                   n@�z�G��?             $@        �       �                   b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     >@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  �H���x�?����C�?M��}t��?e���?��B���?6�����?��RJ)��?���Zk��?;�;��?ى�؉��?�q�q�?�q�q�?      �?                      �?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?�?�?e�kBP��?�	A����?
���F�?��F($�?�������?�������?�q�q�?�q�q�?�m۶m��?�$I�$I�?      �?      �?              �?      �?        ���Kh�?h/�����?��y��y�?�a�a�?      �?                      �?      �?              �?              �?        <<<<<<�?�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��:��:�?_�_��?vb'vb'�?;�;��?      �?      �?              �?��8��8�?�8��8��?�rO#,��?|a���?�5��P�?y�5���?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?]t�E]�?F]t�E�?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��8��8�?�q�q�?      �?              �?      �?      �?              �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?      �?6�d�M6�?e�M6�d�?n۶m۶�?I�$I�$�?�q�q�?9��8���?              �?�������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?l(�����?(������?�������?�?      �?        ى�؉��?;�;��?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?              �?      �?                      �?�c�1Ƹ?�s�9��?�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �$e��?¶��>�?��ۥ���?6��9�?]t�E�?t�E]t�?      �?      �?颋.���?�.�袋�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?vb'vb'�?;�;��?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?۶m۶m�?%I�$I��?�q�q�?9��8���?              �?      �?      �?              �?      �?      �?              �?      �?        (�����?�5��P�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?                      �?      �?        ��L�Ϻ?a�|���?mާ�d�?2�h�>�?�"Qj�a�?��Z9��?              �?[�R�֯�?��+j�?�����?�ȍ�ȍ�?�a�a�?=��<���?UUUUUU�?UUUUUU�?;�;��?;�;��?(�����?�5��P�?              �?      �?      �?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?        �?�?(�����?�5��P�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�?�?      �?      �?              �?      �?                      �?��!XG�?XG��).�?�a�a�?�<��<��?;�;��?ى�؉��?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?��Moz��?��,d!�?      �?        F]t�E�?/�袋.�?�������?�������?              �?      �?      �?              �?      �?      �?              �?      �?              �?        ى�؉��?��؉���?      �?        m�w6�;�?r1����?�������?�������?      �?        �������?�������?333333�?ffffff�?      �?      �?              �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKǅ�h��B�1         B                   �`@�#i����?�           ��@               )                    �?����m�?�            �r@              "                    �Q@�b��gS�?�             m@                                 i@h�WH��?�             k@                                   �?`���i��??             V@       ������������������������       �        1            �Q@               
                    �?�t����?             1@              	                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                  pi@     ��?T             `@        ������������������������       �                     @                                  ``@��U!~2�?R            �^@                                   �?�>4և��?%             L@                                    L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                   @L@H%u��?              I@       ������������������������       �                     <@                                   _@���!pc�?             6@        ������������������������       �                     $@                                   �?      �?	             (@        ������������������������       �                     @        ������������������������       �                     @                                   �?�����?-            �P@        ������������������������       �                      @               !                 ����? ����?,            @P@                                   �l@؇���X�?             @                                    J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        '             M@        #       (                   �i@     ��?
             0@        $       %                    �?�<ݚ�?             "@        ������������������������       �                     �?        &       '                   �_@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        *       5                 ����?������?.            @Q@       +       4                    `Q@�t����?             A@       ,       3       
             �?�g�y��?             ?@       -       2                    �?�nkK�?             7@        .       /                   �n@ףp=
�?             $@       ������������������������       �                     @        0       1                   Hq@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        6       A       
             �?z�G�z�?            �A@       7       8                    X@��a�n`�?             ?@        ������������������������       �                     �?        9       @                    �?��S�ۿ?             >@        :       ;                    �?"pc�
�?             &@        ������������������������       �                     @        <       ?                    @N@      �?              @        =       >                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                     @        C       �                    �?F�Q�j�?           {@       D       �                 ���@��:x���?�            �r@       E       x       
             �?��򟜠�?�            Pq@       F       q                    �?�+$�jP�?t            �g@       G       n                    �?Xf`�>��?b            �d@       H       m                   �f@���(\��?`             d@       I       J                    �?      �?X             b@        ������������������������       �                     D@        K       f       	             �?D>�Q�?A             Z@        L       _                 ����?�	j*D�?              J@       M       X                    @L@�7����?            �G@       N       W                    �?6YE�t�?            �@@       O       V                    �?д>��C�?             =@       P       U                    �?`2U0*��?             9@       Q       T                    @D@���7�?             6@        R       S                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        Y       ^                    �?և���X�?             ,@       Z       [                    �?���Q��?             $@        ������������������������       �                      @        \       ]                   �b@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        `       a                   �`@���Q��?             @        ������������������������       �                     �?        b       e                   �o@      �?             @       c       d                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        g       h                   �? ��WV�?!             J@       ������������������������       �                    �F@        i       l                   �a@����X�?             @        j       k                   p`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        o       p                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        r       s                    �?� �	��?             9@        ������������������������       �                     $@        t       u                   `\@��S�ۿ?
             .@       ������������������������       �                     &@        v       w                   �l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        y       �                   �c@`���i��?-             V@        z                        ����?�7��?            �C@       {       |                   @[@$�q-�?             :@        ������������������������       �                     �?        }       ~                    a@`2U0*��?             9@       ������������������������       �                     8@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                    �H@        ������������������������       �                     4@        �       �       
             �?��M���?\             a@       �       �                   d@Ʋ(>^�?B            @W@       �       �                    �?HP�s��?4            �R@        �       �                   �b@8�Z$���?             :@       �       �                    �?�����?             5@        ������������������������       �                     @        �       �                 ����?�r����?             .@        �       �                 `ff�?�<ݚ�?             "@       �       �                    �H@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �c@���Q��?             @       �       �                   Po@�q�q�?             @        ������������������������       �                     �?        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?@9G��?             �H@       �       �                   `h@�X�<ݺ?             B@        �       �                   `g@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     <@        ������������������������       �                     *@        �       �                    �?X�<ݚ�?             2@       �       �                   �^@���|���?             &@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @        �       �                   0a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �c@�+��<��?            �E@       �       �                    �M@�n_Y�K�?             :@       �       �                    �?z�G�z�?	             .@        ������������������������       �                     @        �       �                    �?�z�G��?             $@       �       �                     H@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���|���?             &@       �       �                    �?���Q��?             $@        ������������������������       �                     @        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 hff @@�0�!��?             1@       �       �                    �?@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        �       �                   Pd@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�b��"     h�h)h,K ��h.��R�(KK�KK��hi�Bp  �5�;���?%e��?��JH7�?M�I�-2�?����˽?�i��F�?B{	�%��?��^B{	�?F]t�E�?F]t�E�?              �?�?<<<<<<�?�q�q�?9��8���?              �?      �?                      �?      �?     ��?      �?        鰑�?����-��?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?        ���Q��?)\���(�?              �?t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?���@��?g��1��?      �?         �����? �����?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?9��8���?�q�q�?              �?      �?      �?      �?                      �?              �??���(�?ہ�v`��?<<<<<<�?�?��{���?�B!��?�Mozӛ�?d!Y�B�?�������?�������?      �?              �?      �?              �?      �?              �?              �?                      �?�������?�������?�c�1Ƹ?�s�9��?      �?        �?�������?F]t�E�?/�袋.�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        H��c���?q�*8���?1ogH���?;Cb�ΐ�?��� ù�?��M���?/�����?B{	�%��?�cp>��?dp>�c�?ffffff�?�����̼?      �?      �?      �?        b'vb'v�?vb'vb'�?vb'vb'�?;�;��?]AL� &�?G}g����?'�l��&�?e�M6�d�?a���{�?|a���?���Q��?{�G�z�?�.�袋�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?      �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?              �?      �?      �?                      �?              �?�������?333333�?      �?              �?      �?      �?      �?      �?                      �?              �?O��N���?;�;��?      �?        �m۶m��?�$I�$I�?      �?      �?              �?      �?              �?              �?              �?      �?              �?      �?        )\���(�?�Q����?      �?        �?�������?              �?      �?      �?      �?                      �?F]t�E�?F]t�E�?��[��[�?�A�A�?�؉�؉�?;�;��?              �?���Q��?{�G�z�?      �?                      �?      �?              �?                      �?�������?�?EM4�D�?/���.�?{�G�z�?q=
ףp�?;�;��?;�;��?�a�a�?=��<���?              �?�?�������?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?9/���?������?�q�q�?��8��8�?      �?      �?              �?      �?                      �?              �?�q�q�?r�q��?F]t�E�?]t�E]�?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?w�qG��?w�qG�?ى�؉��?;�;��?�������?�������?              �?333333�?ffffff�?      �?      �?      �?                      �?      �?      �?      �?                      �?]t�E]�?F]t�E�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ZZZZZZ�?�������?n۶m۶�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK݅�h��B@7         �                    �?"��G,�?�           ��@                                 �g@�*�@P��?            {@               
                    �?�Km�a̾?T            �a@                                   �?���|���?             &@                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     @               	                   Pe@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?���f�?L             `@                                  �?�eGk�T�?8            �W@                                  �b@ ���J��?            �C@       ������������������������       �                     A@                                  �Y@z�G�z�?             @        ������������������������       �                      @                                   �?�q�q�?             @                     
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        !             L@                                  c@�t����?             A@                                 �]@`Jj��?             ?@       ������������������������       �        
             1@                      	             �?؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @                                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                �                    �?d}h���?�            `r@       !       D                    �?��u���?�            Pq@        "       )                   pi@.}Z*�?/            �Q@        #       $       
             �?      �?              @        ������������������������       �                     @        %       (                    �?z�G�z�?             @       &       '                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        *       1                    �?���h%��?*            �O@        +       0                    �?؇���X�?
             ,@        ,       /                 @33�?      �?             @       -       .                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        2       C                    �?ZՏ�m|�?             �H@       3       4                 ����?������?             A@        ������������������������       �                     @        5       B                    @P@����X�?             <@       6       A                    �?�ՙ/�?             5@       7       @                   0o@D�n�3�?             3@       8       ;                    �?�q�q�?
             (@       9       :                    �K@      �?              @        ������������������������       �                      @        ������������������������       �                     @        <       =                    �G@      �?             @        ������������������������       �                     �?        >       ?                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@        E       x                   �a@=�Ѝ;�?u            �i@       F       G                   �Q@���*�?H             ^@        ������������������������       �                      @        H       I                    Z@�:�B��?G            �]@        ������������������������       �        	             1@        J       w                    �?@�G��S�?>            @Y@       K       n                    �?�GN�z�?7             V@       L       M                     H@��oh���?*            @R@        ������������������������       �        
             2@        N       Y                    _@�1�`jg�?             �K@        O       T                    p@��S���?             .@       P       S                   �k@�z�G��?             $@        Q       R                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        U       V                    �?z�G�z�?             @        ������������������������       �                      @        W       X                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       k                    �?R���Q�?             D@       [       `                   `a@l��
I��?             ;@        \       _                    `@8�Z$���?             *@        ]       ^                    �M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        a       b                    �?և���X�?	             ,@        ������������������������       �                      @        c       j                    �?      �?             (@       d       e                    ]@�eP*L��?             &@        ������������������������       �                     @        f       g                    �?����X�?             @        ������������������������       �                     �?        h       i                    �L@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        l       m                   �q@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        o       p                   �a@������?             .@       ������������������������       �                     "@        q       r                 ����?�q�q�?             @        ������������������������       �                     @        s       t                    �?�q�q�?             @        ������������������������       �                     �?        u       v                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        y       �                    �? �#�Ѵ�?-            �U@       z       �                   pl@$Q�q�?"            �O@        {       �                    �?"pc�
�?             6@       |       }                   �b@������?	             1@        ������������������������       �                     @        ~       �                    �?�	j*D�?             *@               �                    �?և���X�?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �D@        ������������������������       �                     7@        �       �                    �?j���� �?
             1@        ������������������������       �                     @        �       �                    �?      �?             ,@        ������������������������       �                     @        �       �                 ����?      �?              @        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    I@DE��2{�?�            �r@        �       �       	             �?؇���X�?            �A@       �       �                   @b@     ��?             @@       �       �                    �Q@`Jj��?             ?@       �       �                 `ff�?(;L]n�?             >@       ������������������������       �                     6@        �       �                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 Zff�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @L@��%p���?�            �p@       �       �                    �? �M*k�?~            �h@       �       �                   �g@p�`Bh�?a            �b@       �       �       
             �?p���?`            �b@       ������������������������       �        :            �V@        �       �                   0n@����˵�?&            �M@       ������������������������       �                     >@        �       �                   �[@ܷ��?��?             =@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        ������������������������       �                     �?        �       �                    �?��+7��?             G@        ������������������������       �                     "@        �       �                   l@4�B��?            �B@        �       �                    �?�n_Y�K�?             *@       �       �                   �g@�q�q�?             (@        ������������������������       �                     @        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                   0k@r�q��?             @        ������������������������       �                     @        �       �                    @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             8@       �       �                    �?�X�<ݺ?             2@       ������������������������       �        
             *@        �       �                   0q@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                    �H@���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?�������?'             Q@       �       �                   �?`��}3��?            �J@       �       �                    b@���N8�?             E@       �       �                   �_@�r����?             >@        �       �                   �^@�z�G��?             $@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        �       �                    `P@      �?             (@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                   ht@��S�ۿ?
             .@       ������������������������       �                     (@        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  �UK���?U�)|��?��Tx*<�?���a���?PuPu�?_�_��?F]t�E�?]t�E]�?      �?      �?              �?      �?        �������?�������?              �?      �?        ��=aOأ?�'�	{��?�X�0Ҏ�?��=�ĩ�?�A�A�?��-��-�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�?<<<<<<�?�B!��?���{��?              �?�$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?I�$I�$�?�A��}�?���ޓ��?�
��V�?�z2~���?      �?      �?      �?        �������?�������?      �?      �?      �?                      �?      �?        EQEQ�?v]�u]��?۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        9/����?�>4և��?�?xxxxxx�?              �?�$I�$I�?�m۶m��?�a�a�?�<��<��?(������?l(�����?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?              �?R�yY�'�?������?wwwwww�?""""""�?      �?        �pR���?�c+����?              �?z��~�X�?�Q`ҩ�?]t�E�?�袋.��?����?ȏ?~��?              �?��)A��?��k߰�?�������?�?333333�?ffffff�?333333�?�������?              �?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?h/�����?Lh/����?;�;��?;�;��?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?      �?t�E]t�?]t�E�?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?                      �?;�;��?�؉�؉�?              �?      �?        �?wwwwww�?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?�}A_Ч?�/����?AA�?~��}���?F]t�E�?/�袋.�?�?xxxxxx�?              �?;�;��?vb'vb'�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?              �?�������?ZZZZZZ�?      �?              �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ,�Œ_,�?O贁N�?�$I�$I�?۶m۶m�?      �?      �?�B!��?���{��?�?�������?              �?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?$�q���?q��;2l�?J�f�?n�%��ʴ?���M�&�?ـl@6 �?\���(\�?{�G�z�?      �?        W'u_�?��/���?      �?        ��=���?a���{�?      �?      �?              �?      �?              �?                      �?zӛ����?Y�B��?      �?        �Y7�"��?L�Ϻ��?ى�؉��?;�;��?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?UUUUUU�?��8��8�?�q�q�?      �?        �������?�������?      �?                      �?      �?      �?333333�?�������?      �?              �?      �?              �?      �?                      �?�������?�������?�琚`��?M0��>��?�a�a�?��y��y�?�������?�?ffffff�?333333�?      �?              �?      �?      �?                      �?ffffff�?�������?      �?                      �?      �?      �?              �?      �?        F]t�E�?]t�E]�?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��B�;         d                    �?�#i����?�           ��@               9                    �?t�F�}�?�            Pv@                                   �?H}m�y��?W            �a@                                  �q@�E��ӭ�?             B@                                  �?8�Z$���?             :@                                 `Z@      �?
             0@        ������������������������       �                     @                      	             �?$�q-�?	             *@       	       
                   `c@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                   �?���Q��?             $@                                 �r@�q�q�?             "@        ������������������������       �                     @                                  `c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?               ,                   P`@���΍L�?C            �Z@                                 �a@�5��?#             K@        ������������������������       �                     1@                                  Pc@�Gi����?            �B@                      
             �?r�q��?             (@                               033@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               '                   �^@�q�����?             9@              &                   �f@�t����?
             1@               %                    �?؇���X�?	             ,@       !       $                     F@"pc�
�?             &@        "       #                    @B@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        (       )                    �L@      �?              @       ������������������������       �                     @        *       +                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        -       .                   �c@4��?�?              J@       ������������������������       �                     B@        /       4                    �?     ��?	             0@        0       3                   �c@      �?              @       1       2                   �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        5       8                    �?      �?              @        6       7                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        :       Y                    �?�V���?�            �j@       ;       X                 ���@�i�y�?w            �g@       <       Q                    �O@ �%�}��?v            �g@       =       B                   @[@P����?p             f@        >       ?                   �Z@r�q��?             @       ������������������������       �                     @        @       A                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        C       D                    �?�h%�M��?j            `e@        ������������������������       �                      I@        E       N                    �?p�,�V��?J            @^@       F       M                   �a@�6H�Z�?G            @]@        G       H       	             �?�(\����?             D@        ������������������������       �        	             5@        I       L                    �?�}�+r��?             3@       J       K                   pa@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        1            @S@        O       P                 `ff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        R       W                    �?"pc�
�?             &@       S       V                 ����?����X�?             @        T       U                    a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        Z       ]                    `@ȵHPS!�?             :@        [       \       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ^       _                   @f@���7�?             6@       ������������������������       �                     1@        `       a       
             �?z�G�z�?             @        ������������������������       �                     @        b       c                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       �                 ����?�^����?�            �w@        f       w                   a@���0��?I             [@        g       l                   �Z@���!pc�?             F@        h       i                   �[@      �?
             0@       ������������������������       �                     @        j       k                    @L@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        m       v                    �?؇���X�?             <@        n       u                    �O@      �?              @       o       p                    �?z�G�z�?             @        ������������������������       �                      @        q       r                 ����?�q�q�?             @        ������������������������       �                     �?        s       t                   `X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        x       �                   �b@     8�?*             P@        y       z                   `Y@ףp=
�?             >@        ������������������������       �                     �?        {       �                   @s@ 	��p�?             =@       |       }                     M@h�����?             <@       ������������������������       �                     9@        ~                           �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?��.k���?             A@        �       �                    �?�����H�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             9@        �       �                   �b@�����H�?             "@       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?     ��?             0@       �       �                   �`@��
ц��?
             *@        �       �                    �?      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ]@r�q��?             @        ������������������������       �                     @        �       �                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�Jx���?�            �p@        �       �                    �?���N8�?             E@       �       �                   `^@؇���X�?            �A@        �       �                    �?      �?             @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   hs@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   pc@ 	��p�?             =@       �       �                 033�? 7���B�?             ;@        ������������������������       �                     (@        �       �                    �?��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        �       �                   `t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `T@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    ]@�K�w���?�            `l@        �       �                     H@tk~X��?             B@        �       �                    �?��
ц��?             *@       �       �                    �?�<ݚ�?             "@       �       �                    \@      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    Y@�nkK�?             7@       ������������������������       �        	             ,@        �       �                   @Z@�����H�?             "@        ������������������������       �                     @        �       �                   �k@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pe@ �r�ɻ?{            �g@       �       �                    �?�tVV�?y            �g@       �       �                   �Q@��AV���?k            �d@        �       �                   Pa@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@���ׇD�?i            �d@       �       �                 ����?pY���D�?f            �c@        �       �                    �L@���Q��?             @        ������������������������       �                     �?        �       �                   �i@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@`#`��k�?a             c@       �       �                    �?�x�E~�?8            @V@       ������������������������       �        .            �R@        �       �                    �?�r����?
             .@       �       �                   �\@؇���X�?	             ,@        �       �                   @V@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �        )             P@        �       �                   pd@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pm@؇���X�?             5@       �       �                    S@�KM�]�?             3@       �       �                    �L@r�q��?             (@       ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  �5�;���?%e��?777777�?�������?e�v�'��?΁D+l�?�q�q�?r�q��?;�;��?;�;��?      �?      �?              �?�؉�؉�?;�;��?      �?      �?      �?                      �?      �?              �?        �������?333333�?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?                      �?      �?        ��sHM�?�	�[��?/�����?h/�����?              �?o0E>��?#�u�)��?�������?UUUUUU�?�m۶m��?�$I�$I�?      �?                      �?      �?        ���Q��?�p=
ף�?�������?�������?�$I�$I�?۶m۶m�?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ى�؉��?�N��N��?              �?      �?      �?      �?      �?�������?�������?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?D��=��?��V!�n�?�������?AA�?]AL� &�?m�w6�;�?�V'u�?'u_[�?�������?UUUUUU�?      �?              �?      �?      �?                      �?��/��?@��?      �?        ˠT�x�?���k��?�������?���?333333�?�������?      �?        �5��P�?(�����?�؉�؉�?;�;��?      �?                      �?      �?              �?              �?      �?              �?      �?        /�袋.�?F]t�E�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?��N��N�?�؉�؉�?      �?      �?      �?                      �?�.�袋�?F]t�E�?      �?        �������?�������?      �?              �?      �?      �?                      �?�X%�,.�?é��t��?����K�?���Kh�?t�E]t�?F]t�E�?      �?      �?              �?�q�q�?�q�q�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?     ��?      �?�������?�������?              �?������?�{a���?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?      �?�؉�؉�?�;�;�?      �?      �?      �?      �?      �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �f�P���?'s�M��?��y��y�?�a�a�?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?�{a���?������?h/�����?	�%����?              �?�?�������?              �?      �?              �?      �?              �?      �?        �m۶m��?�$I�$I�?              �?      �?        ����L�?�hAjv�?9��8���?r�q��?�؉�؉�?�;�;�?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        d!Y�B�?�Mozӛ�?              �?�q�q�?�q�q�?              �?UUUUUU�?�������?      �?                      �?o��2�|�?�ќ5(�?br1���?ڨ�l�w�?7Āt,e�?��8���?UUUUUU�?UUUUUU�?      �?                      �?8��18�?�cp>�?�3���?a~W��0�?�������?333333�?      �?              �?      �?              �?      �?        p�pŊ?@�?��?p�\��?����G�?              �?�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?UUUUUU�?�������?      �?                      �?�$I�$I�?۶m۶m�?(�����?�k(���?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK�h��B�<         �                    �?�#i����?�           ��@                                 @E@<=�h)W�?           �{@                                   �?z�G�z�?'            @P@                                   �?���>4��?             <@                                  �?������?
             1@              	                    �?      �?	             0@                                 �d@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        
                           �?�q�q�?             @                                 `Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                    �B@               g                 pff�?B��u��?�            �w@              4                    �?t�l�ϡ�?�            �r@                                  @j@�d�K���?(            �P@                                  @\@b�2�tk�?             2@        ������������������������       �                     @                                ����?������?
             .@                                  c@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                  �b@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @               /                    �?�J��%�?            �H@              &                   xp@���N8�?             E@               #       	             �?ȵHPS!�?             :@       !       "                    @F@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �        
             6@        $       %                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        '       (                   a@     ��?
             0@        ������������������������       �                     @        )       *                    �?���|���?             &@        ������������������������       �                     @        +       ,                   Hq@�q�q�?             @        ������������������������       �                     �?        -       .                    f@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        0       1                   �`@؇���X�?             @        ������������������������       �                     @        2       3                 @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        5       X                    @M@�|����?�            `m@       6       S       	             �?8��$��?z            �g@       7       >                   0n@�>����?A             [@       8       =       
             �?@	tbA@�?(            @Q@        9       <                   �\@ ��WV�?             :@        :       ;                   g@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             4@        ������������������������       �                    �E@        ?       R                    �?:�&���?            �C@       @       I                    �?tk~X��?             B@       A       H                   0c@PN��T'�?             ;@        B       G                    �?���|���?             &@        C       F                 ����?�q�q�?             @       D       E                   �[@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        J       M                    @F@�q�q�?             "@        K       L                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        N       Q                    �?r�q��?             @       O       P                    �L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       U                   �?��'�`�?9            �T@       ������������������������       �        6            �S@        V       W                   0p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        Y       ^                   Pc@���!pc�?             F@       Z       ]                   `_@`2U0*��?             9@        [       \                   �n@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        _       f                 033�?D�n�3�?	             3@       `       e                    �?ҳ�wY;�?             1@       a       d                   0d@և���X�?             ,@       b       c                   �Z@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        h       }                    �?\I�~�?1            @S@       i       l                    �?��V�I��?            �G@        j       k                   `Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        m       |                 ��� @Hث3���?            �C@       n       y                   �n@���@M^�?             ?@       o       x                   @b@��<b���?             7@       p       q                   �]@�t����?             1@        ������������������������       �                      @        r       w                   �`@z�G�z�?             .@       s       v                   �a@؇���X�?             ,@        t       u                   pf@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        z       {                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ~       �                    �?z�G�z�?             >@              �                    �?�����H�?             ;@        �       �                    �?����X�?             @        �       �                 ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?P���Q�?             4@       ������������������������       �                     &@        �       �                 ����?�����H�?             "@        �       �                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����? ]�к��?�             r@        �       �                    �?v�(��O�?)            �R@       �       �                 ����?�3Ea�$�?             G@       �       �                   �b@�X�<ݺ?             B@       ������������������������       �                     A@        ������������������������       �                      @        �       �                    �M@�z�G��?             $@       �       �                    p@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?V�a�� �?             =@        �       �       	             �?���Q��?             $@       �       �                    �?      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�KM�]�?             3@       �       �                   �c@�IєX�?	             1@       ������������������������       �                     &@        �       �                    h@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�'�%c�?�            �j@       �       �                   �b@Ά^���?i            �b@       �       �                    �?�T�H���?_            �`@       �       �                    �N@ȖLy�r�?^            �`@       �       �                    �?�	��)��?G            �Y@        �       �                   �j@��
ц��?
             *@        ������������������������       �                     @        �       �                 ����?���Q��?             $@       �       �                    �?����X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �^@�q�q�?             @        ������������������������       �                     �?        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ����?ףp=
�?=            �V@        �       �                    c@z�G�z�?            �A@       �       �                    �?ܷ��?��?             =@       �       �                    �?�>����?             ;@       ������������������������       �                     1@        �       �                    �?z�G�z�?             $@        �       �                   @_@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @^@h㱪��?$            �K@        �       �                   �\@�t����?
             1@        ������������������������       �                      @        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     C@        ������������������������       �                     ?@        ������������������������       �                     �?        �       �                    �?��S���?
             .@       �       �                   �c@�n_Y�K�?	             *@        �       �                    q@�q�q�?             @       �       �                   �m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �e@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @N@ ����?)            @P@       ������������������������       �                    �C@        �       �                   �`@ ��WV�?             :@       ������������������������       �                     3@        �       �                    �?؇���X�?             @       �       �                    �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  �5�;���?%e��?�I .Ԝ�?el��W��?�������?�������?n۶m۶�?I�$I�$�?xxxxxx�?�?      �?      �?;�;��?;�;��?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?              �?B-'r��?}��U��?L%�S��?�jg����?����?�rv��?�8��8��?9��8���?              �?wwwwww�?�?      �?      �?              �?      �?        /�袋.�?F]t�E�?      �?                      �?9/����?c}h���?��y��y�?�a�a�?�؉�؉�?��N��N�?d!Y�B�?�Mozӛ�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        {��#�?�7'�h�?vX�Q�}�?�x��* �?�Kh/��?h/�����?�%~F��?ہ�v`��?O��N���?;�;��?�������?UUUUUU�?              �?      �?              �?              �?        �A�A�?�o��o��?r�q��?9��8���?&���^B�?h/�����?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?              �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?�������?�������?      �?                      �?      �?              �?        1P�M��?��k���?      �?              �?      �?      �?                      �?F]t�E�?t�E]t�?���Q��?{�G�z�?�������?�������?      �?                      �?      �?        (������?l(�����?�������?�������?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?                      �?      �?        �cj`��?!��O���?G}g����?r1����?      �?      �?              �?      �?        ��-��-�?�i�i�?�s�9��?�c�1��?��,d!�?��Moz��?�������?�������?              �?�������?�������?۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?      �?                      �?      �?              �?      �?      �?                      �?              �?�������?�������?�q�q�?�q�q�?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?�������?ffffff�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?        �y�!���?�!����?O贁N�?Y�%�X�?��,d!�?����7��?�q�q�?��8��8�?              �?      �?        ffffff�?333333�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?��{a�?a���{�?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �k(���?(�����?�?�?      �?        �������?UUUUUU�?              �?      �?              �?      �?      �?                      �?X:Ɂ���?���O�m�?��:m��?K~���?t��:W�?R�ߦ5�?�1���?���-�j�?r^�	��?ch���V�?�؉�؉�?�;�;�?              �?333333�?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �������?�������?�������?�������?a���{�?��=���?h/�����?�Kh/��?              �?�������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��)A��?־a���?�?<<<<<<�?              �?�q�q�?9��8���?              �?      �?                      �?              �?      �?        �������?�?ى�؉��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?         �����? �����?              �?;�;��?O��N���?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         �                    �?�/�$�y�?�           ��@              i       	             �?�|�tr��?	           `z@              6                    �?�S.���?�            �q@               +                 033�?���X�K�?Y            �`@                                  �?>A�F<�?J            �\@                     
             �?Pq�����?7            @U@                                   �M@r�q��?             (@               	                    �?      �?             @        ������������������������       �                     �?        
                          @]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                  �t@��pBI�?0            @R@                                  �?�k~X��?/             R@                                  �^@h�����?             <@                                  `c@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                      F@        ������������������������       �                     �?               *                   �r@�f7�z�?             =@                                  �?�q�q�?             8@                                  m@�C��2(�?	             &@                               `ff�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   _@��
ц��?             *@        ������������������������       �                      @                )       
             �?���|���?             &@       !       "                   b@X�<ݚ�?             "@        ������������������������       �                     @        #       (                    �?�q�q�?             @       $       %                    �L@z�G�z�?             @        ������������������������       �                     @        &       '                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ,       5                 ���
@؇���X�?             5@       -       4                   @b@ףp=
�?             4@       .       /                   �d@�}�+r��?             3@       ������������������������       �        	             .@        0       3                   ``@      �?             @        1       2                     I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        7       \                    �? �T�7��?_            �b@       8       E                    �?6�iL�?I            �]@       9       D                   0a@���Lͩ�?+            �R@       :       ;                   �h@��0{9�?             �G@        ������������������������       �                     6@        <       =                 ����? �o_��?             9@       ������������������������       �        
             ,@        >       C                 ����?���|���?	             &@       ?       B                   �_@      �?              @        @       A                 @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     <@        F       [                    �?�K��&�?            �E@       G       P                    �?      �?             D@       H       O                    `P@�GN�z�?             6@       I       L                 hff�?�KM�]�?             3@       J       K                   pf@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        M       N                   0l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Q       Z                 033�?X�<ݚ�?             2@       R       U                    �?      �?
             0@        S       T                    @M@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        V       Y                   `m@z�G�z�?             $@        W       X                    @F@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ]       d                    �?     ��?             @@        ^       c                   �e@@�0�!��?             1@        _       b                    ^@      �?             @       `       a                 @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        e       f                    l@��S�ۿ?             .@       ������������������������       �        	             (@        g       h                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        j       u                    �?�u����?Q             a@       k       t                   @g@���͡?C            @\@       l       m                    �?����X�?B             \@        ������������������������       �                     :@        n       o                    @L@��f�{��?2            �U@       ������������������������       �        /            �T@        p       s                    q@      �?             @       q       r                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        v                           �?r�q��?             8@       w       x                   �W@ҳ�wY;�?	             1@        ������������������������       �                     @        y       ~                   �c@      �?             (@       z       }                   �^@�q�q�?             "@        {       |                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �M@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �D@:ө�!��?�            �s@        �       �                    @C@ҳ�wY;�?	             1@        ������������������������       �                     @        �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �W@�a�3u>�?�            pr@        ������������������������       �                      @        �       �                    �?�6hܟo�?�            Pr@        �       �                    �?���|���?             F@       �       �                    �J@"pc�
�?            �@@        �       �                   �`@�q�q�?             (@        �       �                    k@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �`@���N8�?             5@        �       �                     N@r�q��?             @       ������������������������       �                     @        �       �                   `^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             .@        �       �                    �?�C��2(�?             &@       ������������������������       �                     "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?н����?�             o@       �       �                    �R@��$xtW�?�            �j@       �       �                    a@P�S�L�?�            `j@       �       �                    _@p��ճC�?n             f@        �       �                   �o@�ʈD��?            �E@       �       �                   �g@�g�y��?             ?@       ������������������������       �                     6@        �       �                    �?�����H�?             "@        ������������������������       �                     �?        �       �                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �J@      �?             (@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �s@@M^l���?W            �`@       ������������������������       �        Q            @_@        �       �       
             �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   po@b�h�d.�?            �A@       �       �                   �m@���!pc�?             6@       �       �                   @b@�S����?             3@       �       �                    �?      �?
             0@        ������������������������       �                      @        ������������������������       �        	             ,@        �       �                    \@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                      @        �       �                   �\@*O���?             B@        ������������������������       �                     @        �       �       
             �?*;L]n�?             >@       �       �                    �?��}*_��?             ;@       �       �                   @b@և���X�?             5@       �       �                    �?�t����?             1@        ������������������������       �                     @        �       �                   pf@؇���X�?
             ,@       �       �                    _@$�q-�?	             *@        �       �                    ]@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                 `ff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�Bp  L�f���?Z�L��?��p�C�?�Tx��?� �6_�?4�i�A��?l�l��?�'}�'}�?������?Cy�5��?~~~~~~�?�?�������?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ���Ǐ�?����?�8��8��?�q�q�?�m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?                      �?a���{�?O#,�4��?�������?�������?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?�؉�؉�?�;�;�?      �?        F]t�E�?]t�E]�?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?�������?�������?(�����?�5��P�?              �?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        t�@��?�Œ_,��?'u_[�?ylE�pR�?�K~��?�6�i�?L� &W�?m�w6�;�?              �?�Q����?
ףp=
�?              �?]t�E]�?F]t�E�?      �?      �?      �?      �?              �?      �?              �?                      �?              �?��)kʚ�?���)k��?      �?      �?�袋.��?]t�E�?�k(���?(�����?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?r�q��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?      �?                      �?      �?      �?ZZZZZZ�?�������?      �?      �?      �?      �?      �?                      �?              �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        <�H��?"��uy�?$��Co�?x�!���?n۶m۶�?�$I�$I�?      �?        ������?�}A_Ї?      �?              �?      �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?i�i��?��[��[�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?���5n�?C��r$:�?      �?        �L��Y�?���Z�i�?F]t�E�?]t�E]�?F]t�E�?/�袋.�?�������?�������?      �?      �?              �?      �?              �?      �?              �?      �?        �a�a�?��y��y�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?]t�E�?F]t�E�?      �?              �?      �?      �?                      �?�����?�a�E���?��n�?�?����?JQ/#��?`�
��T�?]t�E�?]t�E�?�}A_з?A_���?�B!��?��{���?              �?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?      �?333333�?�������?      �?                      �?              �?����~?&���g��?              �?      �?      �?              �?      �?        _�_��?;��:���?t�E]t�?F]t�E�?^Cy�5�?(������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �q�q�?�q�q�?              �?�������?""""""�?B{	�%��?_B{	�%�?۶m۶m�?�$I�$I�?�������?�������?      �?        �$I�$I�?۶m۶m�?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?              �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKυ�h��B�3         z                    �?���
%�?�           ��@              m       	             �? ��7E��?           �z@              "                    �?P����?�            y@                                  �`@�y(dD�?'            @P@                                   �?��>4և�?             <@                     
             �?��+7��?             7@                                 �R@և���X�?
             ,@        ������������������������       �                     @        	       
                    �?���!pc�?             &@        ������������������������       �                     �?                                   �?�z�G��?             $@        ������������������������       �                     @                                   �I@և���X�?             @                               ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @                                   @G@�MI8d�?            �B@        ������������������������       �                      @                      
             �?(N:!���?            �A@                               ���@XB���?             =@       ������������������������       �        
             1@                                  �\@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@               !                    �?      �?             @                                  Pd@      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        #       Z                    �?ؙ/,T�?�             u@       $       9                    �?@����<�?�            �q@        %       .                    �G@��a��?O            @^@        &       '                     E@և���X�?             @        ������������������������       �                      @        (       -                    �?���Q��?             @       )       *                    �?      �?             @        ������������������������       �                     �?        +       ,                   (p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        /       6                 033@P�Lt�<�?J            �\@       0       5                   �^@�K}��?A            �Y@        1       4                   �h@@4և���?	             ,@        2       3                     N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        8             V@        7       8                   @U@r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        :       O       
             �?�Q��k�?e             d@       ;       <                    @K@0�ޤ��?S            @`@       ������������������������       �        +             P@        =       D                    �?���7�?(            �P@        >       C                    �?؇���X�?	             ,@       ?       @                 ����?"pc�
�?             &@        ������������������������       �                     @        A       B                   �\@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        E       N                    �? pƵHP�?             J@       F       M                    �?��Y��]�?            �D@       G       L                    �M@�(\����?             D@        H       I                    @M@P���Q�?             4@       ������������������������       �        	             1@        J       K                    a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                     &@        P       Y                 `ff�?�r����?             >@       Q       X                   c@���|���?
             &@       R       S                   `]@X�<ݚ�?             "@        ������������������������       �                     @        T       W                    @K@�q�q�?             @       U       V                   �r@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        [       \                    S@t�6Z���?!            �K@        ������������������������       �                     �?        ]       d                    �?H�ՠ&��?              K@        ^       c                    �?�n_Y�K�?	             *@       _       b                    �P@      �?              @       `       a                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        e       l                    �R@������?            �D@       f       g                   @a@�(\����?             D@       ������������������������       �                    �A@        h       k                    �?z�G�z�?             @       i       j                 033@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        n       u                   �`@      �?             >@       o       p                   @]@�<ݚ�?
             2@        ������������������������       �                     @        q       r                    �L@��S�ۿ?             .@       ������������������������       �                     &@        s       t                   @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        v       y                     K@�8��8��?             (@        w       x                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        {       �                    �?�˱��H�?�            �r@       |       �                    �?��k�c��?�            `o@       }       �                    @M@����p�?�            �i@       ~       �                    �?`�g����?o             f@              �                   @[@0�`G�r�?e            `d@        �       �       	             �?8�Z$���?	             *@       �       �                    �?      �?              @       �       �                    �F@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@p���?\            �b@       �       �                   �b@`����֜?V            �a@       �       �                    @ 
�V�?Q            �`@       ������������������������       �        P            �`@        ������������������������       �                     �?        �       �                   �f@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �_@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?8�Z$���?
             *@       ������������������������       �                     $@        �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@����X�?             <@        �       �                    �?��
ц��?             *@        ������������������������       �                     @        �       �                 ����?���Q��?             $@       �       �                    �N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����?�r����?             .@       �       �       
             �?�8��8��?             (@       ������������������������       �                     "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    q@��|�5��?!            �G@       �       �                    \@ܷ��?��?             =@        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    @I@�q�q�?             @        ������������������������       �                     �?        �       �                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �e@ �q�q�?             8@       ������������������������       �                     .@        �       �       
             �?�����H�?             "@       ������������������������       �                     @        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �r@X�<ݚ�?	             2@       �       �       
             �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?
j*D>�?             J@       �       �                    @N@�\��N��?             C@       �       �                   `_@X�Cc�?             <@        ������������������������       �                     *@        �       �       
             �?�q�q�?	             .@       �       �                   �b@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                   `a@؇���X�?	             ,@       ������������������������       �                     &@        �       �                    _@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��\���?��Q���?:�����?q����?����i��?J���h�?Wj�Vj��?�J��J��?۶m۶m�?I�$I�$�?zӛ����?Y�B��?�$I�$I�?۶m۶m�?              �?F]t�E�?t�E]t�?      �?        ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?�������?333333�?      �?                      �?      �?              �?                      �?L�Ϻ��?��L���?      �?        �A�A�?|�W|�W�?�{a���?GX�i���?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?      �?      �?              �?      �?              �?                      �?1�0ð?z��y���?��|G��?3��g�?���|���?��2(&�?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?(�����?���k(�?�?�������?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?              �?UUUUUU�?�������?      �?                      �?ffffff�?�������?z�z��?/�B/�B�?              �?F]t�E�?�.�袋�?�$I�$I�?۶m۶m�?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?              �?      �?                      �?;�;��?'vb'vb�?������?8��18�?�������?333333�?�������?ffffff�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?�?�������?F]t�E�?]t�E]�?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?��)A��?X���oX�?      �?        {	�%���?������?ى�؉��?;�;��?      �?      �?�������?UUUUUU�?      �?                      �?              �?              �?������?p>�cp�?�������?333333�?              �?�������?�������?      �?      �?      �?                      �?              �?      �?              �?      �?9��8���?�q�q�?              �?�������?�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?l����?O���!��?oI�!m��?���򖄺?�������?�����Ҳ?�袋.��?]t�E]�?*�/��?�E:i�?;�;��?;�;��?      �?      �?333333�?�������?      �?                      �?      �?              �?        \���(\�?{�G�z�?�������?�A�A�?������?g��1�~?      �?                      �?�������?UUUUUU�?      �?                      �?�������?�������?              �?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?�;�;�?�؉�؉�?      �?        �������?333333�?�������?�������?              �?      �?                      �?�������?�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?br1���?x6�;��?��=���?a���{�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?UUUUUU�?      �?        �q�q�?�q�q�?      �?              �?      �?      �?                      �?r�q��?�q�q�?�������?�������?              �?      �?              �?        ;�;��?b'vb'v�?y�5���?�5��P�?%I�$I��?�m۶m��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?              �?        �������?�������?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKㅔh��B�8         d                    �?�r,��?�           ��@                                  �^@�8~��?�            t@               
       
             �?��R[s�?            �A@                                   �?�n_Y�K�?             *@                                  �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?               	                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?"pc�
�?             6@                                433�?���!pc�?             &@                                   �?      �?             @        ������������������������       �                     �?                                   п�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  p`@�C��2(�?             &@       ������������������������       �                     "@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               ;                 pff�?&�cm���?�            �q@              4                    �?L���
B�?�            �i@              '                    �?�+?�?~            �g@                                   �?����X�?             <@                                   �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?               "       
             �?     ��?
             0@                !                    �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        #       $                    �?r�q��?             @       ������������������������       �                     @        %       &                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       1                   �t@@3����?m            @d@       )       0                    �?�Fǌ��?j            �c@        *       -                    �? ��WV�?"             J@       +       ,                   �f@@��8��?             H@       ������������������������       �                    �G@        ������������������������       �                     �?        .       /                   ``@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        H            �Z@        2       3                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        5       6                    ]@�t����?             1@        ������������������������       �                     @        7       :                 ����?�eP*L��?             &@       8       9                    �?X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        <       K                    �?V�K/��?4            �S@        =       D       
             �?R�}e�.�?             :@        >       C                   �o@�eP*L��?             &@       ?       B                    �?X�<ݚ�?             "@       @       A                   �e@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        E       F                    �?��S�ۿ?	             .@       ������������������������       �                     "@        G       J                    �?r�q��?             @        H       I                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        L       ]       	             �?r�z-��?#            �J@       M       R                    �?      �?             @@        N       Q                 ����?����X�?             @        O       P                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        S       \                   �s@ �o_��?             9@       T       W                    �?��<b���?             7@       U       V                   �b@�S����?             3@       ������������������������       �                     0@        ������������������������       �                     @        X       [                    �?      �?             @       Y       Z                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ^       c                    �?����X�?             5@       _       b                    �L@ҳ�wY;�?
             1@       `       a                    @      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        e       �                    �??d)�?�            �y@        f       �                 ����?�,����?W             b@        g       z                   d@�ګH9�?+            �Q@       h       y                    �?H%u��?             I@       i       j                    �?=QcG��?            �G@        ������������������������       �                     "@        k       p                    �?�˹�m��?             C@       l       o                   �b@���}<S�?             7@       m       n                    `P@���7�?             6@       ������������������������       �        
             5@        ������������������������       �                     �?        ������������������������       �                     �?        q       x                 ����?��S�ۿ?	             .@       r       s                   �`@@4և���?             ,@        ������������������������       �                      @        t       u                    �?r�q��?             @        ������������������������       �                     @        v       w                     P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        {       |                 `ffֿև���X�?             5@        ������������������������       �                      @        }       �                   �b@�\��N��?             3@       ~                           \@���Q��?
             .@        ������������������������       �                     �?        �       �                   �q@X�Cc�?	             ,@       �       �                    b@�<ݚ�?             "@       �       �                    �?      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   0a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��G���?,            �R@       �       �                   @u@f.i��n�?            �F@       �       �                    �O@R���Q�?             D@       �       �                    @     ��?             @@       �       �                    b@�û��|�?             7@       �       �                   �_@�E��ӭ�?             2@       �       �                    @J@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                    �?�q�q�?             @       �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    S@z�G�z�?             @        ������������������������       �                      @        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     =@        �       �                    �?�NJa&��?�            �p@        �       �                   �R@>��C��?            �E@        ������������������������       �                     @        �       �                   `a@�d�����?             C@        �       �                   a@���Q��?             4@        �       �                   �`@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?8�Z$���?             *@       �       �                    �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                 ����?�����H�?             2@       �       �                    �H@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��S�ۿ?�             l@        �       �                 ����?8�Z$���?&            @P@        ������������������������       �                     >@        �       �                    �?����X�?            �A@        �       �                    �?@4և���?
             ,@       ������������������������       �                     "@        �       �                   �h@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    b@և���X�?             5@       ������������������������       �                     &@        �       �                 ����?ףp=
�?             $@        �       �                    @M@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@      �?d             d@       �       �                    �? ���v��?>            �X@       �       �                   �j@�(\����?2             T@        �       �                   `_@������?            �D@       ������������������������       �                     6@        �       �                    �K@�KM�]�?
             3@       �       �                   �i@�X�<ݺ?	             2@       ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                 033�?�S����?             3@        �       �                    �H@���Q��?             @        ������������������������       �                     �?        �       �                    `@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@4և���?             ,@       �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        &            �N@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  �292ȯ�?�f����?�(��L��?����f��?PuPu�?X|�W|��?ى�؉��?;�;��?�$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?/�袋.�?t�E]t�?F]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?��p���?k��<B��?��pK͆�?�{��ɳ?\���%�?Fڱa��?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�������?�������?      �?                      �?UUUUUU�?�������?              �?      �?      �?              �?      �?        ���Kh�?h/�����?1���M��?�3���?O��N���?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?              �?              �?      �?      �?                      �?�������?�������?      �?        t�E]t�?]t�E�?�q�q�?r�q��?              �?      �?              �?        �Z܄��?�ґ=�?'vb'vb�?�;�;�?]t�E�?t�E]t�?r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�?      �?        �������?UUUUUU�?      �?      �?              �?      �?              �?        �琚`��?����!�?      �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        �Q����?
ףp=
�?��Moz��?��,d!�?^Cy�5�?(������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �$I�$I�?�m۶m��?�������?�������?      �?      �?      �?                      �?              �?              �?L	e�h��?����%��?�(ٵ���?�k%�6�?e�v�'��?6��9�?)\���(�?���Q��?x6�;��?AL� &W�?      �?        ��P^Cy�?^Cy�5�?ӛ���7�?d!Y�B�?�.�袋�?F]t�E�?      �?                      �?              �?�������?�?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?              �?�5��P�?y�5���?333333�?�������?              �?%I�$I��?�m۶m��?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?333333�?              �?      �?                      �?v�)�Y7�?#�u�)��?�>�>��?�`�`�?�������?�������?      �?      �?��,d!�?8��Moz�?r�q��?�q�q�?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?                      �?IT�n�?~5&��?qG�w��?$�;��?              �?y�5���?Cy�5��?�������?333333�?۶m۶m�?�$I�$I�?      �?                      �?;�;��?;�;��?UUUUUU�?�������?      �?                      �?              �?�q�q�?�q�q�?�������?�������?      �?        �q�q�?�q�q�?              �?      �?      �?              �?      �?                      �?�?�������?;�;��?;�;��?              �?�$I�$I�?�m۶m��?�$I�$I�?n۶m۶�?              �?�������?�������?              �?      �?        ۶m۶m�?�$I�$I�?              �?�������?�������?�������?�������?      �?                      �?      �?              �?      �?1ogH�۩?�y;Cb�?�������?333333�?������?p>�cp�?              �?(�����?�k(���?�q�q�?��8��8�?              �?      �?              �?                      �?^Cy�5�?(������?�������?333333�?      �?              �?      �?              �?      �?        �$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B@.                             �?T8���?�           ��@                                   �?�<ݚ��?_             b@                               ���@pY���D�?6            �S@       ������������������������       �        4            @S@        ������������������������       �                      @                                  �b@� ���?)            @P@                                  �?�t����?            �I@              	                   @[@��|�5��?            �G@        ������������������������       �                      @        
                           @D@z�G�z�?            �F@        ������������������������       �                     �?                      	             �?"pc�
�?             F@                                 `a@�<ݚ�?             B@                                  �?H%u��?             9@       ������������������������       �                     (@                                  �a@�θ�?             *@        ������������������������       �                     "@                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?�eP*L��?             &@                               ����?؇���X�?             @                                 Hr@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             ,@               h                    �?2� J��?p           p�@               W                   �b@�qu}+�?�            �v@       !       8                   P`@��ӿ���?�            �s@       "       +                    �?p�����?�             n@        #       $                   �_@�8��8��?&             N@        ������������������������       �                     <@        %       &                 ����?     ��?             @@       ������������������������       �                     7@        '       *                    �?X�<ݚ�?             "@       (       )                   �p@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ,       7                    �?�o"Q9a�?q            �f@        -       0                 `ff�? >�֕�?            �A@        .       /                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                   �[@Pa�	�?            �@@        ������������������������       �                     1@        3       4                    �R@      �?	             0@       ������������������������       �                     (@        5       6       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        ^            @b@        9       <                   �`@h�˹�?2             S@        :       ;                   �`@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        =       V       
             �?$�q-�?,            @P@       >       C                    �?`�H�/��?%            �I@        ?       B                    ^@      �?             @        @       A                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        D       U                    @M@dP-���?!            �G@       E       R                    @L@�����H�?             B@       F       M                    �?��S�ۿ?             >@       G       L                   �a@ 7���B�?             ;@       H       I                 033�?��S�ۿ?             .@        ������������������������       �                     @        J       K                   �m@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        N       O                    Z@�q�q�?             @        ������������������������       �                     �?        P       Q                   (p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       T                 hff�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     ,@        X       ]                 hff�?X��ʑ��?            �E@        Y       Z                   �d@z�G�z�?             .@       ������������������������       �                     $@        [       \                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ^       c                    j@��X��?             <@        _       b                    �?����X�?             @        `       a                    W@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        d       e                   �`@��s����?             5@       ������������������������       �                     .@        f       g                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        i       �                   @E@�����?�            �l@        j              	             �?�!���?             A@       k       ~                    �O@r֛w���?             ?@       l       u                 ����?V�a�� �?             =@        m       n                    @D@X�<ݚ�?             "@        ������������������������       �                      @        o       t                    �J@և���X�?             @       p       q                     G@z�G�z�?             @        ������������������������       �                     �?        r       s                   Pa@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        v       w                    �?ףp=
�?             4@        ������������������������       �                     &@        x       }                    �?�<ݚ�?             "@        y       z                    �M@�q�q�?             @        ������������������������       �                     �?        {       |                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?y            �h@        �       �       	             �?�1�`jg�?$            �K@       �       �                    �?�99lMt�?            �C@       �       �                   �c@�LQ�1	�?             7@       �       �                 833@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �?     ��?             0@       �       �                    �?      �?             $@       �       �                   �f@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �H@      �?             0@       ������������������������       �                     "@        �       �                    f@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?dP-���?U            �a@       �       �                   �f@��b�h8�?L            �_@       �       �                 ���@�.ߴ#�?I            �^@       �       �                   Pd@(;L]n�?H             ^@       �       �                    �?P���Q�?.             T@       �       �                    _@(�5�f��?-            �S@        �       �                   �a@HP�s��?             9@        �       �       	             �?�<ݚ�?             "@       ������������������������       �                     @        �       �                   �^@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             0@        �       �       
             �?@3����?             K@       ������������������������       �                    �A@        �       �                   �c@�}�+r��?             3@       ������������������������       �                     0@        �       �                 `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     D@        ������������������������       �                      @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	             �?����X�?	             ,@       �       �                    �?���|���?             &@       �       �                 033�?      �?              @       �       �                   �d@�q�q�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  6n����?�� ���?�q�q�?�8��8��?a~W��0�?�3���?      �?                      �?�����?�ȍ�ȍ�?�������?�������?br1���?x6�;��?              �?�������?�������?              �?/�袋.�?F]t�E�?9��8���?�q�q�?)\���(�?���Q��?      �?        ى�؉��?�؉�؉�?      �?              �?      �?              �?      �?        t�E]t�?]t�E�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?                      �?              �?�|����?��w�;�?[�[��?�I��I��?-hk�ש?}I��b�?$�$��?���?UUUUUU�?UUUUUU�?              �?      �?      �?              �?r�q��?�q�q�?�m۶m��?�$I�$I�?      �?                      �?              �?�rS�<��?6��{��?�A�A�?��+��+�?      �?      �?              �?      �?        |���?|���?              �?      �?      �?              �?      �?      �?      �?                      �?              �?�5��P�?^Cy�5�?F]t�E�?]t�E]�?              �?      �?        ;�;��?�؉�؉�?�?�������?      �?      �?      �?      �?      �?                      �?              �?W�+�ɵ?�����F�?�q�q�?�q�q�?�?�������?h/�����?	�%����?�?�������?              �?�q�q�?�q�q�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�}A_�?��}A�?�������?�������?              �?333333�?�������?      �?                      �?n۶m۶�?%I�$I��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?z��y���?�a�a�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�@�V���?�����a�?�������?�������?�B!��?���{��?a���{�?��{a�?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?�������?�������?      �?              �?      �?      �?                      �?              �?�������?�������?              �?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?        ۶m۶m�?�$I�$I�?��k߰�?��)A��?5H�4H��?�o��o��?��Moz��?Y�B��?��y��y�?�a�a�?      �?                      �?              �?      �?      �?      �?      �?UUUUUU�?�������?              �?      �?              �?                      �?      �?      �?      �?        �m۶m��?�$I�$I�?      �?                      �?�����F�?W�+�ɵ?������?�@ �?�K�`m�?XG��).�?�������?�?ffffff�?�������?�=Q���?�&��jq�?q=
ףp�?{�G�z�?9��8���?�q�q�?      �?        333333�?�������?      �?                      �?      �?        ���Kh�?h/�����?      �?        �5��P�?(�����?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?333333�?�������?      �?                      �?�m۶m��?�$I�$I�?]t�E]�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         �       
             �?�[��N�?�           ��@                                  �?�"�&z�?`           8�@                                   �?���5��?c            �c@                                 �g@��(\���?M             ^@                               pff�?�1e�3��?L            �]@       ������������������������       �        >            @Y@                                   @M@j���� �?             1@              	                    �?�����H�?             "@        ������������������������       �                     @        
                           �?z�G�z�?             @                                  �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                  �^@<ݚ)�?             B@        ������������������������       �                     &@                                   �O@� �	��?             9@                                 �p@�t����?             1@                                  �?X�<ݚ�?             "@                                  �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                   `@      �?              @        ������������������������       �                      @        ������������������������       �                     @                U                    �?��t���?�            �x@        !       D                    @N@ޚ)�?^             b@       "       /                   �a@
j*D>�?D             Z@        #       (                    Z@�C��2(�?            �@@        $       '                    �?����X�?             @        %       &                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        )       .                 ����? ��WV�?             :@       *       +                    �?�8��8��?
             (@       ������������������������       �                     "@        ,       -                   Pa@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        0       =                    �?L�];�?.            �Q@       1       :                   �r@�����?             E@       2       7                   �e@ >�֕�?            �A@       3       6                    f@Pa�	�?            �@@        4       5                   @_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        8       9                   @m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ;       <                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        >       ?                    �?ܷ��?��?             =@       ������������������������       �                     7@        @       C                    �?      �?             @        A       B                    @L@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        E       R                   0c@R���Q�?             D@       F       O                    �?������?            �B@       G       H                   `]@l��\��?             A@        ������������������������       �        
             1@        I       N                    �?@�0�!��?             1@       J       M                   �m@և���X�?             @       K       L                 ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        P       Q                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        S       T                 033@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        V       g                    �?X����?�            `o@        W       f                    �?д>��C�?$             M@       X       Y                    `@�4�����?             ?@        ������������������������       �                     (@        Z       [                    �?�\��N��?             3@        ������������������������       �                     @        \       a                    �?     ��?             0@        ]       `                    �?և���X�?             @       ^       _                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        b       e                    @K@X�<ݚ�?             "@       c       d                    b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        h       �                   ``@�-j'�?{             h@        i       t                    �?h�V���?8             V@        j       m                    �?�z�G��?             $@        k       l                   @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        n       o                 ����?�q�q�?             @        ������������������������       �                     �?        p       q                 ����?z�G�z�?             @        ������������������������       �                     @        r       s                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       �                    �?$�q-�?1            �S@       v                          0i@��ɉ�?(            @P@        w       ~                    �?���}<S�?             7@       x       }                    \@      �?             0@        y       |                   @`@����X�?             @       z       {                   �^@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     E@        �       �                 ���@�	j*D�?	             *@       �       �                    �?"pc�
�?             &@       �       �                   �[@�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �K@      �?              @        ������������������������       �                     @        �       �                   �X@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?@��!�Q�?C            @Z@       �       �                   �a@�\=lf�?.            �P@        �       �                    �?`2U0*��?             9@        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   �h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     E@        ������������������������       �                     C@        �       �                    @L@dP,k|��?g            �f@       �       �                    �?��E��?@            �\@       �       �                 ����?$�q-�?-            �V@       �       �                    �?��
���?'            �R@       �       �                    @G@      �?              P@        ������������������������       �                    �@@        �       �                    �?`Jj��?             ?@        ������������������������       �                     $@        �       �                    �G@�����?             5@        ������������������������       �                      @        ������������������������       �        
             3@        ������������������������       �                     &@        �       �                    �?     ��?             0@        ������������������������       �                     "@        �       �                    V@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 @33�?8����?             7@        ������������������������       �                     @        �       �                   P`@j���� �?             1@        �       �                 ����?      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             "@        �       �                   �b@\X��t�?'            @Q@       �       �                 pff�?����X�?            �H@       �       �                    n@�f7�z�?             =@       �       �                 ����?���!pc�?             6@       �       �                    �?z�G�z�?             4@       �       �                    �?������?	             1@       ������������������������       �                     &@        �       �                   �]@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    \@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 033�?ףp=
�?	             4@       �       �                    �?z�G�z�?             $@       �       �                   @e@r�q��?             @       �       �                   p`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   ``@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 ��� @z�G�z�?             4@       �       �                   �a@      �?
             0@        �       �                    `@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�b�      h�h)h,K ��h.��R�(KK�KK��hi�BP  B~�9�J�?�@c�Z�?_� M�?P���o��?i�i��?\��[���?�������?333333�?�/���?W'u_�?      �?        �������?ZZZZZZ�?�q�q�?�q�q�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?              �?�8��8��?��8��8�?              �?)\���(�?�Q����?�������?�������?r�q��?�q�q�?�������?UUUUUU�?      �?                      �?              �?              �?      �?      �?              �?      �?        ^-n����?�td�@T�?��8��8�?9��8���?;�;��?b'vb'v�?F]t�E�?]t�E�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?;�;��?O��N���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?SO�o�z�?Zas �
�?=��<���?�a�a�?��+��+�?�A�A�?|���?|���?�������?�������?              �?      �?              �?              �?      �?              �?      �?        �m۶m��?�$I�$I�?      �?                      �?a���{�?��=���?              �?      �?      �?      �?      �?      �?                      �?              �?333333�?333333�?к����?��g�`��?�������?------�?              �?�������?ZZZZZZ�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?���e�?�_FA@s�?|a���?a���{�?��RJ)��?���Zk��?              �?y�5���?�5��P�?      �?              �?      �?۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?              �?�q�q�?r�q��?UUUUUU�?�������?              �?      �?              �?                      �?�1�K��?��LF�W�?/�袋.�?�袋.��?333333�?ffffff�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�? �����??�?��?d!Y�B�?ӛ���7�?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?              �?              �?              �?;�;��?vb'vb'�?F]t�E�?/�袋.�?�q�q�?9��8���?      �?              �?      �?              �?      �?      �?      �?                      �?              �?      �?        8�8��? �����?g��1��?"=P9���?{�G�z�?���Q��?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?��|�(�?��ݮ�?���b:��?1��t��?�؉�؉�?;�;��?&�X�%�?O贁N�?      �?      �?      �?        ���{��?�B!��?      �?        =��<���?�a�a�?              �?      �?              �?              �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?        8��Moz�?d!Y�B�?              �?ZZZZZZ�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?��Moz��?!Y�B�?�$I�$I�?�m۶m��?a���{�?O#,�4��?t�E]t�?F]t�E�?�������?�������?�?xxxxxx�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �������?�������?�������?�������?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?      �?              �?      �?                      �?�������?�������?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�}�JhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK텔h��B@;         r                    �?�_y���?�           ��@              e                    �?^��4m�?�             w@                                  �?h
WY�v�?�            �s@               	                    T@�ƫ�%�?:            @V@                                  @b@z�G�z�?             @                                 �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        
                           �M@ ��N8�?7             U@       ������������������������       �        /             R@                                   �?�8��8��?             (@        ������������������������       �                     @                                  �c@z�G�z�?             @        ������������������������       �                     @                                  �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               T                    �?�����?�            �l@              S                   �g@������?~             i@              :                    @L@(1�Fh�?}            �h@                                  �?D��*�4�?Z            @a@                     	             �?@uvI��?=            �X@                                  pf@�?�|�?            �B@       ������������������������       �                     ;@                                  `]@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        '            �N@               -                    �?R���Q�?             D@               (                    @F@      �?             4@                !                    @D@և���X�?             @        ������������������������       �                     �?        "       %                    @E@      �?             @        #       $                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        &       '                   `i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        )       ,                    �?$�q-�?             *@       *       +                    T@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        .       7                   �e@z�G�z�?             4@       /       2                   @_@�t����?             1@        0       1                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       6                    �?��S�ۿ?             .@       4       5                    �?@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?        ������������������������       �                     �?        8       9                    �D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ;       L                    �?����S��?#             M@       <       E       	             �?�����?             C@       =       D                   p@����X�?             <@       >       C                   �`@z�G�z�?             9@        ?       B                   �a@X�<ݚ�?             "@       @       A                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     @        F       I                   Hp@���Q��?             $@       G       H                     Q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        J       K                    q@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        M       P                   �n@      �?             4@       N       O                    e@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        Q       R                   p`@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        U       V                    �?��S���?             >@        ������������������������       �                     $@        W       ^                   (p@z�G�z�?             4@       X       [                    �?؇���X�?
             ,@       Y       Z                   �d@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        \       ]                    @M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        _       d                 ����?�q�q�?             @        `       a                    �?�q�q�?             @        ������������������������       �                     �?        b       c                    �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        f       o                    �R@>a�����?!            �I@       g       n                    �?�q��/��?             G@        h       i                   �f@X�<ݚ�?             "@        ������������������������       �                     @        j       m                    �?r�q��?             @       k       l                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �B@        p       q                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        s       �                   �b@؇���X�?�            �v@       t       �                    �?�1h�'��?�            `r@       u       �                 ����?���H��?�            @j@       v       {                   0f@r�q��?^            @a@        w       x       
             �?(;L]n�?             >@       ������������������������       �                     :@        y       z                   @e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        |       �                   Pi@�{��?��?G             [@        }       ~                    �D@�	j*D�?
             *@        ������������������������       �                      @               �                   @_@"pc�
�?             &@        �       �                   @`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?\�ih�<�?=            �W@        �       �                   (s@�q�q�?             8@       �       �       	             �?z�G�z�?             4@       �       �                   �`@�S����?             3@        �       �                   �l@      �?             @        ������������������������       �                     �?        �       �                   �\@���Q��?             @        ������������������������       �                     �?        �       �                    [@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        �       �                   �v@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @K@@�j;��?,            �Q@        �       �                    n@Pa�	�?            �@@        �       �                   �\@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     4@        �       �                   �a@�?�'�@�?             C@       �       �                    �?������?            �B@        ������������������������       �                      @        �       �       	             �?\-��p�?             =@       �       �                   �[@؇���X�?             <@        �       �       
             �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����?���N8�?             5@        �       �                 `ff�?؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   b@������?,             R@       ������������������������       �        %             P@        �       �                   �b@      �?              @       �       �                    �?���Q��?             @       �       �                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? ��N8�?2             U@        �       �                    n@�IєX�?             1@       ������������������������       �        
             (@        �       �                    �M@z�G�z�?             @        ������������������������       �                     @        �       �                   (p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        $            �P@        �       �                   0c@<=�,S��?+            �Q@        �       �                    `@      �?              @        �       �                    @B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   X~@V��z4�?&             O@       �       �                     P@��0u���?%             N@       �       �                    �?J��D��?"             K@        �       �       
             �?�E��ӭ�?             2@       �       �                    @K@�θ�?             *@        �       �                    �D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    b@�����H�?             "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �_@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     K@�q�q�?             B@       �       �                     E@r�q��?             2@       �       �       
             �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?      �?
             2@       �       �                   `d@�	j*D�?             *@       �       �                   d@      �?              @       �       �                    �?�q�q�?             @       �       �       	             �?z�G�z�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  V�.�#��?աh6n��?�|����?�S�n�?��f����?�e�}��?��x�3�?�as�ì?�������?�������?      �?      �?              �?      �?                      �?�y��y��?�a�a�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?              �?      �?      �?                      �?�T>��u�?���(�?
ףp=
�?ףp=
��?������?h�����?ہ�v`��?)�3J���?�Cc}h��?9/���?*�Y7�"�?к����?      �?        �������?�������?              �?      �?              �?        �������?�������?      �?      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?      �?              �?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?<<<<<<�?�?      �?      �?      �?                      �?�������?�?n۶m۶�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        X�i���?O#,�4��?Q^Cy��?^Cy�5�?�m۶m��?�$I�$I�?�������?�������?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?333333�?�������?�������?UUUUUU�?      �?                      �?      �?      �?              �?      �?              �?      �?�������?�?      �?                      �?�������?333333�?              �?      �?                      �?�������?�?      �?        �������?�������?�$I�$I�?۶m۶m�?�������?�������?              �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�?�������?��Mozӻ?�B����?r�q��?�q�q�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?333333�?�������?              �?      �?        �$I�$I�?۶m۶m�?�E�_���?K���+�?��y��y�?�0�0�?UUUUUU�?�������?�?�������?              �?      �?      �?              �?      �?        /�����?���^B{�?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?        Ai�
��?�%N���?�������?�������?�������?�������?^Cy�5�?(������?      �?      �?      �?        �������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?              �?      �?      �?                      �?H���@��?w�'�K�?|���?|���?;�;��?�؉�؉�?      �?                      �?              �?y�5���?������?к����?��g�`��?              �?�{a���?a����?�$I�$I�?۶m۶m�?۶m۶m�?�$I�$I�?      �?                      �?�a�a�?��y��y�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?              �?      �?        �q�q�?�q�q�?              �?      �?      �?�������?333333�?      �?      �?      �?                      �?      �?                      �?�a�a�?�y��y��?�?�?              �?�������?�������?              �?      �?      �?      �?                      �?              �?X|�W|��?�A�A�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �s�9��?2�c�1�?""""""�?�������?_B{	�%�?�^B{	��?r�q��?�q�q�?�؉�؉�?ى�؉��?      �?      �?              �?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?              �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?      �?;�;��?vb'vb'�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?              �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ'J�OhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKӅ�h��B�4         P                 ����?<���m�?�           ��@               5                    �?V7�`A�?�            �u@              2                   h@��<VO�?�            `o@              +                    �?���C���?�             o@                                  �?���l��?�            �k@                                 @[@p�`Bh�?`            �b@                                  �Z@�θ�?             *@       ������������������������       �                     "@        	       
                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �?�Ŗ�Pw�?X            @a@       ������������������������       �        T            �`@                                  @a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?�ˡ�5��?*            �Q@                                  �?��ϭ�*�?"             M@                                  b@�����H�?            �F@                                  �?������?            �D@       ������������������������       �                     <@                                  �c@8�Z$���?             *@        ������������������������       �                     �?                                   @F@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                  hv@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@               *                    �?��
ц��?             *@               )                 ����?���|���?             &@       !       (                    d@���Q��?             $@       "       '                    �?؇���X�?             @       #       $                   @`@z�G�z�?             @        ������������������������       �                      @        %       &                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ,       1       
             �?���B���?             :@       -       .                    _@     ��?
             0@        ������������������������       �                      @        /       0                     F@d}h���?	             ,@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     $@        3       4                   pn@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        6       ?                    @G@�*v��?>            @X@        7       8                    @D@>���Rp�?             =@        ������������������������       �                     $@        9       :                    �?p�ݯ��?             3@        ������������������������       �                     @        ;       >                    �D@$�q-�?	             *@        <       =       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        @       G                   �a@l��\��?+             Q@       A       B                   �o@p���?             I@       ������������������������       �                     F@        C       D                    �M@r�q��?             @        ������������������������       �                     @        E       F                    `P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        H       O                    �?�E��ӭ�?             2@       I       N       	             �?X�Cc�?             ,@       J       K                    @J@      �?	             (@       ������������������������       �                      @        L       M                    `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        Q       �                    �?�|�+�p�?�             x@        R       w                   �b@�d�K���?\            �`@       S       f                    @M@�G�z.�?7             T@        T       [                 ����?h+�v:�?             A@        U       Z                   @e@r�q��?
             (@       V       Y                   �_@�C��2(�?	             &@        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        \       a                    m@��2(&�?             6@       ]       `                   �^@�X�<ݺ?             2@        ^       _                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        b       e       	             �?      �?             @       c       d                     G@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        g       n                    �?�LQ�1	�?             G@        h       i                   `Z@և���X�?             @        ������������������������       �                     �?        j       m                   �`@�q�q�?             @       k       l                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        o       t       
             �?�7��?            �C@       p       q                    �?(;L]n�?             >@       ������������������������       �                     5@        r       s                 033�?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        u       v                 ����?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        x       �                    �?����0�?%             K@       y       �                    @X�<ݚ�?             B@       z       }                   �d@�+e�X�?             9@       {       |                   Pg@      �?             0@        ������������������������       �                     �?        ������������������������       �        
             .@        ~                           �?X�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @        �       �                   �n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?���Q��?             @       �       �                   @f@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�C��2(�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �e@r�q��?             2@       �       �                    �L@      �?
             0@       ������������������������       �                     *@        �       �                   �e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �U@4�Ջ�;�?�            �o@        ������������������������       �                     �?        �       �                    �? �_�x�?�            `o@        �       �       
             �?�d�����?             C@       �       �                    �?�<ݚ�?             B@        ������������������������       �                     @        �       �                   �a@6YE�t�?            �@@       �       �                   �`@���N8�?             5@       �       �                    �?�n_Y�K�?             *@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@       �       �                   �t@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                      @        �       �                    �?����Q8�?�            �j@       �       �                    �?@9G��?            �h@        �       �                   �b@�����H�?             B@       �       �                   P`@Pa�	�?            �@@        �       �                   �\@      �?              @        ������������������������       �                     @        �       �                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     9@        ������������������������       �                     @        �       �                   i@�(\����?i             d@        ������������������������       �        #            �M@        �       �                    b@��'cy�?F            @Y@       �       �                   �[@`Ql�R�??            �W@        �       �                    �K@�8��8��?             (@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pa@����ȫ�?7            �T@        ������������������������       �                    �D@        �       �                 ����?��Y��]�?            �D@        ������������������������       �                     �?        ������������������������       �                     D@        �       �                     N@����X�?             @       �       �                   �b@���Q��?             @        ������������������������       �                     �?        �       �                    �L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?������?             1@        ������������������������       �                     �?        �       �                   �^@     ��?
             0@        �       �                    [@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �_@�8��8��?             (@       ������������������������       �                     @        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  ���>��?�,@��"�? ��2)�?��:����?�Tw�V�?�ZEtJu�?J)��RJ�?���Zk��?��蕱�?5'��Ps�?���M�&�?ـl@6 �?ى�؉��?�؉�؉�?      �?              �?      �?      �?                      �?��?���?ہ�v`�}?      �?        �������?�������?      �?                      �?�RO�o��?H���@��?����=�?|a���?�q�q�?�q�q�?p>�cp�?������?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?        �؉�؉�?�;�;�?F]t�E�?]t�E]�?�������?333333�?�$I�$I�?۶m۶m�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?        ��؉���?ى�؉��?      �?      �?              �?I�$I�$�?۶m۶m�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�i�n�'�?��Id��?GX�i���?�i��F�?              �?Cy�5��?^Cy�5�?      �?        ;�;��?�؉�؉�?      �?      �?              �?      �?                      �?�������?------�?{�G�z�?\���(\�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?r�q��?�q�q�?�m۶m��?%I�$I��?      �?      �?              �?      �?      �?              �?      �?              �?                      �?&��+���?6�5؝�?����?�rv��?ffffff�?ffffff�?xxxxxx�?�������?�������?UUUUUU�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?t�E]t�?��.���?�q�q�?��8��8�?�������?�������?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        Y�B��?��Moz��?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?�A�A�?��[��[�?�?�������?              �?�q�q�?�q�q�?      �?                      �?�q�q�?�q�q�?      �?                      �?�Kh/���?Lh/����?r�q��?�q�q�?R���Q�?���Q��?      �?      �?              �?      �?        �q�q�?r�q��?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�u]�u]�?EQEQ�?      �?        ����0p�?g��1�?y�5���?Cy�5��?�q�q�?9��8���?      �?        e�M6�d�?'�l��&�?��y��y�?�a�a�?ى�؉��?;�;��?              �?r�q��?�q�q�?�������?UUUUUU�?      �?                      �?              �?              �?              �?      �?        ��Vج?O�o�z2�?9/���?������?�q�q�?�q�q�?|���?|���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?333333�?              �?��be�F�?`ҩy���?W�+�ɕ?}g���Q�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?              �?������?������?              �?������?8��18�?      �?                      �?�$I�$I�?�m۶m��?�������?333333�?      �?              �?      �?              �?      �?                      �?�?xxxxxx�?      �?              �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW�ehG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�-         �       	             �?�$���?�           ��@              �       
             �?A��s��?q           �@              N                    �?08`���?            {@                                   �?�������?j            �d@                                   �R@�LQ�1	�?             G@                                  �?�C��2(�?             F@                                 �U@�t����?             A@        ������������������������       �                      @        	       
                    @O@      �?             @@       ������������������������       �                     2@                                  �^@؇���X�?             ,@                                  0o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @               9                 ����?2��(���?N            �]@                                  �a@p�}�ޤ�?2            @R@                                 @E@���H��?             E@                                   �?      �?             @                                 `Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �?�}�+r��?             C@                                    M@      �?
             0@       ������������������������       �                     &@                                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        !       2                   Pd@`՟�G��?             ?@       "       '                    �?ҳ�wY;�?             1@        #       $                    �?      �?             @        ������������������������       �                     �?        %       &                    @M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        (       1                   0d@�θ�?	             *@       )       ,                    �?�z�G��?             $@        *       +                   ``@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        -       0                    �?���Q��?             @       .       /                   `Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        3       8                   �f@d}h���?             ,@       4       7                   �e@�q�q�?             "@       5       6                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        :       ?                    �?*
;&���?             G@        ;       <                    �?���Q��?             @        ������������������������       �                      @        =       >                 `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        @       A                   �`@������?            �D@        ������������������������       �                     6@        B       G                   `a@���y4F�?             3@        C       F                    �?�q�q�?             @       D       E                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        H       I                   Pm@      �?
             0@       ������������������������       �                     $@        J       M                    �?�q�q�?             @       K       L                   pn@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        O       �                    �?��W[�?�            �p@       P       �                    �Q@pb����?x             g@       Q       �                    �?�1j�P�?v            �f@       R       m                 ����?|�e����?p            `e@        S       T                 833�?$]��<C�?1            �Q@        ������������������������       �                     ?@        U       `                    �?��Q��?             D@       V       [                    �?�	j*D�?             :@        W       Z                    �?���Q��?             $@       X       Y                    @N@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        \       _                    �H@      �?             0@        ]       ^                    �F@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             (@        a       l                   �`@և���X�?	             ,@       b       c                    �?���Q��?             $@        ������������������������       �                     @        d       k                     P@և���X�?             @       e       f                    �?      �?             @        ������������������������       �                     �?        g       h                   �[@�q�q�?             @        ������������������������       �                     �?        i       j                   @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        n       w                    �?` A�c̭??             Y@       o       v                    @J@�}��L�?/            �R@        p       u                 ����?h�����?             <@        q       t                   �h@$�q-�?             *@        r       s                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     .@        ������������������������       �                    �G@        x       {                    �H@HP�s��?             9@        y       z                   h@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        |       �                    @O@���7�?             6@       }       �                    �?�C��2(�?             &@        ~                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     &@        �       �                   �c@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        1            �T@        �       �                    �?�G�"�?^            �a@       �       �                    �?B�����?H             Z@       �       �                     Q@P���Q�?3             T@       �       �                   �c@ ���J��?1            �S@       �       �                   �c@`Ӹ����?            �F@       �       �                    �M@`���i��?             F@       ������������������������       �                     ?@        �       �                    ]@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                      @        �       �                   �h@      �?             8@        ������������������������       �                     @        �       �                    �?��.k���?             1@        ������������������������       �                     @        �       �                    �F@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?����>�?            �B@        �       �                    �?���Q��?             .@        �       �                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �`@���7�?             6@       ������������������������       �                     2@        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�摋���?Z             d@       �       �                 ����?�\=lf�?K            �`@       ������������������������       �        F             `@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �n@�q�q�?             ;@       �       �                    �?�	j*D�?             *@        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  �E$�~V�?�����?�w.��?�!��h��?�%���^�?���Kh�?�YΟ���?�0��?Y�B��?��Moz��?F]t�E�?]t�E�?�?<<<<<<�?      �?              �?      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �Bg�Bg�?�z1�z1�?�z��ի�?�
*T��?�0�0�?��y��y�?      �?      �?      �?      �?              �?      �?                      �?�5��P�?(�����?      �?      �?      �?        333333�?�������?      �?                      �?      �?        �1�c��?�s�9��?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?ى�؉��?333333�?ffffff�?�������?�������?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?        8��Moz�?���,d!�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?������?�|����?              �?(������?6��P^C�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?Q�_T��?�t� ]�?�cxq�?Ë��1�?�8xߺ?������?4��\Fs�?�e4���?�'�K=�?6���?              �?ffffff�?�������?;�;��?vb'vb'�?333333�?�������?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?      �?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?333333�?�������?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?���Q��?
ףp=
�?O贁N�?�_,�Œ�?�$I�$I�?�m۶m��?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?              �?              �?{�G�z�?q=
ףp�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?�.�袋�?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?              �?�������?�������?              �?      �?              �?      �?              �?      �?                      �?�2t�n��?T�"��?vb'vb'�?'vb'vb�?ffffff�?�������?��-��-�?�A�A�??�>��?l�l��?F]t�E�?F]t�E�?      �?        �؉�؉�?;�;��?              �?      �?                      �?      �?                      �?      �?      �?              �?�������?�?      �?        �������?�������?      �?                      �?���L�?�u�)�Y�?333333�?�������?      �?      �?              �?      �?              �?        F]t�E�?�.�袋�?              �?      �?      �?      �?                      �?.>9\�?��6Ϳ?"=P9���?g��1��?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?vb'vb'�?;�;��?      �?      �?      �?                      �?�������?�������?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���zhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK녔h��B�:         h                   �`@&I,|-��?�           ��@                                   �?$6HZl�?�            @u@                      	             �?��i#[�?             E@                                  �?П[;U��?             =@                                  �?8�A�0��?             6@                                  �?�eP*L��?             &@        ������������������������       �                      @                                   �?X�<ݚ�?             "@        	                           �?�q�q�?             @       
                          `X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                    Q@�q�q�?             @                                 �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   �?���!pc�?             &@                                433�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@               C                    �?.�w��K�?�            �r@               *                    �?���Q��?@             Y@               )                 ��� @�Ra����?             F@              &                   �p@z�G�z�?             9@              #                     O@ףp=
�?             4@              "                 ����?�X�<ݺ?             2@                !                    @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        $       %                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        '       (                    �R@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     3@        +       2                 ����?      �?)             L@       ,       -                    �      �?             @@        ������������������������       �                     �?        .       /                   �^@�g�y��?             ?@       ������������������������       �                     2@        0       1                    �?$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        3       B       	             �?�q�q�?             8@       4       ;                    �K@�㙢�c�?             7@        5       :                   �c@      �?             @       6       7                    �?      �?             @        ������������������������       �                      @        8       9                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        <       A                    �?�IєX�?             1@       =       >                    `@��S�ۿ?	             .@       ������������������������       �                     *@        ?       @                 033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        D       K                   �[@��:x�ٳ?z            �h@        E       F                   �c@r�q��?             2@       ������������������������       �                     &@        G       H                    �?և���X�?             @        ������������������������       �                     @        I       J                     O@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        L       c                     Q@������?o            �f@       M       b                    �?�D�e���?f            @e@       N       a                   P`@ȑ����?G            @]@        O       P                    �?HP�s��?             I@        ������������������������       �                     *@        Q       V                    �?������?            �B@        R       S                    �?      �?             @        ������������������������       �                      @        T       U                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        W       ^                    @L@�C��2(�?            �@@       X       ]                   �\@ �q�q�?             8@        Y       Z                    @J@r�q��?             @        ������������������������       �                     @        [       \                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             2@        _       `                   �X@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        )            �P@        ������������������������       �                    �J@        d       e                    �?ףp=
�?	             $@       ������������������������       �                     @        f       g                   P`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        i       �                    �?���,���?�            �x@       j       �                 ���@�%��l �?�            @p@       k       n                    �?h�y���?�             o@        l       m                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        o       �                    @M@�� ^ �?�            @n@       p       �                    �?0?R����?}            �j@       q       v                    �?�+�Y�?\            `c@        r       u       
             �?�7��?            �C@        s       t                   �g@�����H�?             2@       ������������������������       �                     0@        ������������������������       �                      @        ������������������������       �                     5@        w       ~                   @[@XB���?C             ]@        x       y                    �?؇���X�?             ,@       ������������������������       �                     "@        z       }                    �?���Q��?             @       {       |       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @               �                    @L@���J��?<            �Y@       ������������������������       �        7            �W@        �       �                   0b@      �?              @        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 hff�?>���Rp�?!             M@       �       �                    P@t/*�?            �G@        ������������������������       �                     @        �       �                    �D@�Ra����?             F@        ������������������������       �                     @        �       �                   �[@������?            �D@        �       �                   0l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �A@        �       �                   �^@�eP*L��?             &@        ������������������������       �                     @        �       �                    b@      �?              @       �       �                   0l@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �c@8^s]e�?             =@       �       �       
             �?�û��|�?             7@       �       �                   �e@��S���?             .@        ������������������������       �                     @        �       �                   a@�q�q�?
             (@        ������������������������       �                      @        �       �                 ����?z�G�z�?             $@       �       �                    �?����X�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    s@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �f@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        �       �                   `f@�Z4���?P            �`@       �       �                   �b@�[�}r�?O            ``@       �       �                    �?d}h���?(            �Q@        �       �                    �I@D�n�3�?
             3@        ������������������������       �                      @        �       �                 ����?���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �       �                   �m@L紂P�?            �I@       �       �                    �?H�V�e��?             A@       �       �                    �?��Q��?             4@        �       �                    �?և���X�?             @        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �K@�θ�?             *@       �       �                    b@�C��2(�?             &@       �       �                   �`@r�q��?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     1@        �       �                 ����?x>ԛ/��?'            �N@       �       �       	             �?">�֕�?            �A@       �       �                    �?��>4և�?             <@       �       �                   �q@�q�q�?             8@       �       �                    �?$�q-�?             *@       ������������������������       �                     &@        �       �                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �s@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@�	j*D�?             :@        �       �                   @p@�eP*L��?             &@       �       �                    N@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pd@�r����?             .@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                    �?      �?             @        ������������������������       �                      @        �       �                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b�`     h�h)h,K ��h.��R�(KK�KK��hi�B�  �"z?+�?���B`��?�������?�������?�a�a�?�<��<��?�{a���?��=���?/�袋.�?颋.���?t�E]t�?]t�E�?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        t�E]t�?F]t�E�?      �?      �?              �?      �?                      �?      �?              �?        ��c.��?Vg�{��?�������?333333�?]t�E�?]t�E]�?�������?�������?�������?�������?�q�q�?��8��8�?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?333333�?�������?              �?      �?                      �?      �?      �?      �?      �?              �?��{���?�B!��?      �?        �؉�؉�?;�;��?      �?                      �?�������?UUUUUU�?d!Y�B�?�7��Mo�?      �?      �?      �?      �?      �?              �?      �?              �?      �?                      �?�?�?�?�������?              �?      �?      �?              �?      �?                      �?      �?        [�R�֯�?
�����?UUUUUU�?�������?              �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?�q�q�?�q�q�?�???????�?���?��~���?{�G�z�?q=
ףp�?              �?к����?��g�`��?      �?      �?              �?      �?      �?      �?                      �?F]t�E�?]t�E�?UUUUUU�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?9��8���?      �?                      �?              �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        W����?R��3�M�?C/�B/��?�B/�B/�?���{��?!�B�?UUUUUU�?UUUUUU�?      �?                      �?���eP*�?����|��?�J�Q���?ޫ-r�	�?�>.����?�=�ѣ?��[��[�?�A�A�?�q�q�?�q�q�?      �?                      �?      �?        GX�i���?�{a���?۶m۶m�?�$I�$I�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ______�?�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �i��F�?GX�i���?�;����?W�+���?              �?]t�E]�?]t�E�?              �?p>�cp�?������?UUUUUU�?UUUUUU�?              �?      �?              �?        ]t�E�?t�E]t�?      �?              �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?        |a���?	�=����?8��Moz�?��,d!�?�������?�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?�$I�$I�?�m۶m��?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        IT�n��?\�՘H�?ˈ>�:��?�����?۶m۶m�?I�$I�$�?(������?l(�����?              �?F]t�E�?t�E]t�?              �?      �?        �������?�������?ZZZZZZ�?iiiiii�?ffffff�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�؉�؉�?ى�؉��?F]t�E�?]t�E�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?                      �?              �?;ڼOq��?�K�`m�?_�_��?�A�A�?۶m۶m�?I�$I�$�?�������?�������?�؉�؉�?;�;��?      �?              �?      �?              �?      �?        ]t�E�?t�E]t�?              �?      �?                      �?      �?        ;�;��?vb'vb'�?t�E]t�?]t�E�?۶m۶m�?�$I�$I�?              �?      �?                      �?�?�������?�q�q�?9��8���?              �?�������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX^khG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKɅ�h��B@2         X                 ����?j8je3�?�           ��@               K                    �?T�h����?�            �u@              4                    �?&ABD��?�            0r@              	                    I@T��mh��?�             l@                                   `P@�G��l��?             5@                                 �Y@d}h���?             ,@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        
       !                    �?�IєX�?�            �i@                                 `a@��AV���?u            �d@                                 0n@@3����?N             [@       ������������������������       �        -            �O@                                  �?`Ӹ����?!            �F@                                  �?`���i��?              F@        ������������������������       �                     @                                   �? ���J��?            �C@                                 0c@��?^�k�?            �A@                                   �G@@4և���?
             ,@                                  �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                     @        ������������������������       �                     �?                                    N@ ,��-�?'            �M@       ������������������������       �                     E@                                   �N@������?             1@        ������������������������       �                      @                                   �t@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        "       %                   i@�MI8d�?            �B@        #       $                    `@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        &       -                    �L@     ��?             @@       '       ,                    �? ��WV�?             :@       (       )                    @I@�X�<ݺ?             2@       ������������������������       �                     &@        *       +                    d@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        .       3                   �c@�q�q�?             @       /       2                   p`@z�G�z�?             @        0       1                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        5       >                    �?"pc�
�?'            �P@        6       7                    �?�eP*L��?
             &@        ������������������������       �                     @        8       9                   �l@r�q��?             @        ������������������������       �                     @        :       =                    �?�q�q�?             @       ;       <                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ?       D       	             �?lGts��?            �K@       @       A                   �o@���.�6�?             G@       ������������������������       �                    �@@        B       C                    @O@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        E       J                 ����?�q�q�?             "@       F       I                    �?      �?              @       G       H                   �_@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        L       W       	             �?���!pc�?%            �K@       M       P                    �?�LQ�1	�?             G@        N       O                    �?�q�q�?	             (@        ������������������������       �                     @        ������������������������       �                      @        Q       R                    �?�IєX�?             A@       ������������������������       �                     9@        S       V                    �?�<ݚ�?             "@       T       U                   �b@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        Y       v                    �?�.�d��?�            @x@        Z       g                    �?X�<ݚ�?'             K@       [       ^                   �\@     ��?             @@        \       ]                    @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        _       f                    �?\-��p�?             =@       `       a                   0c@�>����?             ;@       ������������������������       �        
             0@        b       c                   �Z@"pc�
�?             &@        ������������������������       �                     �?        d       e                   �u@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        h       k                    �?"pc�
�?             6@        i       j                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       s                   �u@�KM�]�?             3@       m       r                    �?�IєX�?             1@       n       q                 ����?      �?             0@        o       p                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     �?        t       u                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        w       �                    �?ˡ��?�            �t@        x       �                    �?���?:            @V@       y       z                   �V@H.�!���?             I@        ������������������������       �                      @        {       �       	             �?     ��?             H@       |       }                    S@���V��?            �F@        ������������������������       �                      @        ~       �                   �b@X�EQ]N�?            �E@              �                   �r@��p\�?            �D@       �       �                 ����?@-�_ .�?            �B@        �       �                     O@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ;@        �       �                    �?      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?�e����?            �C@       �       �                   �^@     ��?             @@        ������������������������       �                     *@        �       �                   pb@D�n�3�?             3@       �       �                   �U@և���X�?             ,@        ������������������������       �                     @        �       �                   �`@�q�q�?             "@        ������������������������       �                     @        �       �                 ����?���Q��?             @       �       �                    d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                   `e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@���m��?�            �n@       �       �                   �[@���7�?~            �k@        �       �                    b@z�G�z�?             9@       �       �                    �?�LQ�1	�?             7@        ������������������������       �                     &@        �       �                    �K@      �?             (@        ������������������������       �                     @        �       �                 033�?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    f@ ���J��?r            `h@       �       �                    _@���e�?n            �g@        �       �                    �J@ >�֕�?            �A@       �       �       	             �?ףp=
�?             4@       �       �                    @�}�+r��?
             3@       ������������������������       �        	             2@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                    @N@��ꤘ�?Z             c@       ������������������������       �        ?             [@        �       �                    �N@����?�?            �F@        �       �                   �m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     E@        �       �       
             �?����X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    j@�q�����?             9@        ������������������������       �                     $@        �       �                   �l@z�G�z�?	             .@        ������������������������       �                     @        �       �                 033@�z�G��?             $@       �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ���Y��?t�S��?����E�?����t�?x(3���?�����?�gE#��?������?1�0��?��y��y�?I�$I�$�?۶m۶m�?              �?      �?                      �?�?�?��8���?7Āt,e�?���Kh�?h/�����?      �?        ?�>��?l�l��?F]t�E�?F]t�E�?      �?        ��-��-�?�A�A�?_�_��?�A�A�?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?              �?      �?              �?              �?              �?                      �?[4���?'u_[�?      �?        xxxxxx�?�?              �?�������?�?      �?                      �?��L���?L�Ϻ��?�������?333333�?      �?                      �?      �?      �?O��N���?;�;��?��8��8�?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?                      �?F]t�E�?/�袋.�?t�E]t�?]t�E�?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�־a�?�<%�S��?Y�B��?���7���?              �?�؉�؉�?ى�؉��?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?�$I�$I�?�m۶m��?              �?      �?                      �?      �?        t�E]t�?F]t�E�?Y�B��?��Moz��?UUUUUU�?UUUUUU�?      �?                      �?�?�?              �?�q�q�?9��8���?�$I�$I�?�m۶m��?      �?                      �?              �?      �?        :*����?q���
|�?r�q��?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?a����?�{a���?�Kh/��?h/�����?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?                      �?              �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?        (�����?�k(���?�?�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?              �?      �?        �rCH��?B#��-N�?7��Mmj�?e%+Y�J�?)\���(�?�(\����?      �?              �?      �?�>�>��?[�[��?      �?        qG�wĽ?w�qG�?��+Q��?�]�ڕ��?к����?S�n0E�?�������?�������?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�A�A�?�-��-��?      �?      �?              �?l(�����?(������?۶m۶m�?�$I�$I�?              �?UUUUUU�?UUUUUU�?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?򸳄���?�iOd �?F]t�E�?�.�袋�?�������?�������?Y�B��?��Moz��?              �?      �?      �?              �?      �?      �?              �?      �?              �?        �A�A�?��-��-�?AL� &W�?����F}�?�A�A�?��+��+�?�������?�������?(�����?�5��P�?              �?      �?              �?                      �?p�p�z? u�u��?              �?l�l��?��I��I�?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?���Q��?�p=
ף�?              �?�������?�������?      �?        ffffff�?333333�?9��8���?�q�q�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQ��dhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKɅ�h��B@2         V                 ����?��}���?�           ��@                                   �?$f����?�            �u@                                  d@�~6�]�?;            @U@                               ����?�r����?3            �R@       ������������������������       �        $             I@               	                    �?���Q��?             9@                                   �L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        
                            O@�q�q�?             5@                                  b@      �?
             0@        ������������������������       �                     &@                                  �b@���Q��?             @        ������������������������       �                     �?                                   �?      �?             @                     
             �?�q�q�?             @        ������������������������       �                     �?                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �\@z�G�z�?             $@        ������������������������       �                     �?                                   f@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                033�pJQg���?�            �p@        ������������������������       �                      @               G                    �?�C��2(�?�            �p@              6                    �?@Ix�<��?�            �m@               /                    �O@�F�l���?x            �g@       !       "                   @n@p�C��?r            �f@       ������������������������       �        J             ]@        #       .                    �?�FVQ&�?(            �P@       $       %                     G@P�2E��?'            @P@        ������������������������       �                     =@        &       -                   0c@�8��8��?             B@        '       (                   �\@z�G�z�?             .@        ������������������������       �                      @        )       *                   �?$�q-�?
             *@       ������������������������       �                     $@        +       ,                    �M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                     �?        0       5                    r@X�<ݚ�?             "@       1       4       	             �?r�q��?             @       2       3                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        7       B                    �?�q��/��?             G@       8       9                    �?��(\���?             D@        ������������������������       �                     @        :       ;                    �?�C��2(�?            �@@        ������������������������       �                      @        <       A                   �b@H%u��?             9@       =       @                    �M@�8��8��?             8@       >       ?                 433�?�nkK�?             7@       ������������������������       �                     6@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        C       F                 @33�?�q�q�?             @       D       E                   �h@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        H       U                   Pd@�5��?             ;@       I       T       
             �?D�n�3�?             3@       J       S                 ����?     ��?             0@       K       P                    �?�q�q�?	             (@       L       O                   �c@      �?              @       M       N                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        Q       R                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        W       �                    a@��(R�?�            �w@       X       e                    �?�J��?�            �l@        Y       `                    �?�f7�z�?             =@       Z       [                   @k@X�Cc�?	             ,@        ������������������������       �                     @        \       _                    �?����X�?             @       ]       ^                    �M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        a       d                   �r@z�G�z�?             .@       b       c                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        f       i                    �?p���?{             i@        g       h                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        j       w                    �?����e��?y            �h@        k       t                    �Q@ >�֕�?            �A@       l       m       
             �?      �?             @@        ������������������������       �                      @        n       s                    �? �q�q�?             8@        o       r                    �?      �?              @        p       q                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        u       v                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        x                           �?������?d            `d@        y       z                     O@P���Q�?             4@       ������������������������       �        	             &@        {       ~                    �?�����H�?             "@       |       }                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        T            �a@        �       �       
             �?i����?[            @c@       �       �       	             �?H�tL��?F            @^@       �       �                    �?Nṧ'
�?8            �W@       �       �                   �a@��<b���?*            @Q@        �       �                    �?���|���?             6@        �       �                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �J@������?
             1@       �       �                    �?X�<ݚ�?             "@        �       �                   Pm@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @I@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@��0{9�?            �G@       �       �                   �g@�'�`d�?            �@@        ������������������������       �                     @        �       �                   �d@R�}e�.�?             :@       �       �                    �?b�2�tk�?             2@       �       �                    \@     ��?	             0@        �       �                    �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    q@�θ�?             *@       ������������������������       �                     @        �       �                    c@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        �       �                   @b@��
ц��?             :@       �       �                    @K@�q�q�?             5@       �       �                   �e@��S���?             .@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pl@���B���?             :@        ������������������������       �                     (@        �       �                 `ff�?X�Cc�?             ,@        �       �                   �e@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                      @        �       �                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 033�?���|���?            �@@        �       �                    �?�IєX�?
             1@       ������������������������       �                     &@        �       �                   �b@r�q��?             @        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   ``@     ��?             0@       �       �                   �_@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  q��H��?��>���?Xx�Wx��?Q�P��?�?999999�?�?�������?              �?�������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?�������?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?        �������?�������?              �?�q�q�?�q�q�?              �?      �?        ���7G��?\�qA��?              �?]t�E�?F]t�E�?(�X�>�?���v��?L�:,��?:kP<�q�?��K��K�?h�h��?      �?        >����?|���?_�^��?z�z��?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?r�q��?�q�q�?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�B����?��Mozӻ?�������?333333�?      �?        ]t�E�?F]t�E�?      �?        )\���(�?���Q��?UUUUUU�?UUUUUU�?�Mozӛ�?d!Y�B�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?h/�����?/�����?(������?l(�����?      �?      �?�������?�������?      �?      �?�������?�������?              �?      �?                      �?      �?      �?              �?      �?                      �?      �?              �?        ��Eh�?{�����?t�?;��?�����?a���{�?O#,�4��?%I�$I��?�m۶m��?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?;�;��?�؉�؉�?      �?                      �?      �?        {�G�z�?\���(\�?      �?      �?      �?                      �?|���?�>����?�A�A�?��+��+�?      �?      �?              �?UUUUUU�?�������?      �?      �?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        )��I� y?<^l	���?�������?ffffff�?              �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?�����?<�����?���!pc�?�
�GN�?#�X�0�?|n�S���?��Moz��?��,d!�?F]t�E�?]t�E]�?�������?�������?              �?      �?        �?xxxxxx�?�q�q�?r�q��?      �?      �?              �?      �?        �������?�������?              �?      �?                      �?L� &W�?m�w6�;�?'�l��&�?6�d�M6�?              �?�;�;�?'vb'vb�?9��8���?�8��8��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?ى�؉��?              �?      �?      �?              �?      �?              �?                      �?              �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?�������?�?      �?      �?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��؉���?ى�؉��?      �?        %I�$I��?�m۶m��?۶m۶m�?�$I�$I�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?        ]t�E]�?F]t�E�?�?�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���lhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK兔h��B@9         j                    �?&I,|-��?�           ��@              M                 ����?���5���?�            �v@                                 @E@Ԯ�̭~�?�             r@                                   �?\X��t�?             7@                                   �?      �?	             (@        ������������������������       �                     @                                   @D@�q�q�?             "@        ������������������������       �                     �?        	       
                    �      �?              @        ������������������������       �                     �?                                   �?؇���X�?             @       ������������������������       �                     @                                   \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �]@�C��2(�?	             &@                                    M@      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               L                   �g@�^;\��?�            �p@              )                    \@�>K�
}�?�            �p@               (                     N@�I�w�"�?             C@                                 �Z@��hJ,�?             A@        ������������������������       �                     &@               '                    @H@��<b���?             7@                                  �?�q�q�?
             (@        ������������������������       �                      @               &                    �?      �?             $@               %                 ����?����X�?             @       !       $                   �c@�q�q�?             @        "       #       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        *       G                    �?�07�r��?�            `l@       +       2                   Hp@��+��?�            �i@       ,       -                    @M@��V9��?c            �a@       ������������������������       �        R            @^@        .       /                    c@ףp=
�?             4@       ������������������������       �                     ,@        0       1                   �i@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        3       4                   �^@�C��2(�?+            �P@        ������������������������       �                     3@        5       6                   `p@��E�B��?             �G@        ������������������������       �                     @        7       8                    �L@t��ճC�?             F@       ������������������������       �                     <@        9       F       	             �?     ��?
             0@       :       E                    �?�z�G��?	             $@       ;       <                   `_@      �?              @        ������������������������       �                     �?        =       B                    �?����X�?             @       >       A       
             �?z�G�z�?             @        ?       @                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        C       D                   @t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        H       I                   `c@      �?             4@        ������������������������       �                     "@        J       K                   Pd@�eP*L��?	             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        N       U                    �?p�ݯ��?0             S@        O       R                   �b@�S����?             C@       P       Q                   �e@�FVQ&�?            �@@       ������������������������       �                     ?@        ������������������������       �                      @        S       T                     P@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        V       [                    �?D�n�3�?             C@        W       X                    �?؇���X�?             @       ������������������������       �                     @        Y       Z                    �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        \       i                 033@�g�y��?             ?@       ]       f                    �?�5��?             ;@       ^       _                    �?@�0�!��?             1@       ������������������������       �                     &@        `       e                 ����?      �?             @       a       d                    �?      �?             @       b       c                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        g       h                    b@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        k       �                   �b@t����?�             w@       l       �                   �a@�F�j��?�            �r@       m       �                    �P@�cX1!��?�             o@       n       �                 ����?`�q��־?�             m@       o       z                    �?�C��2(�?d            @c@        p       y       
             �?�q�q�?
             (@       q       r                   �\@      �?             $@        ������������������������       �                     @        s       x                    @O@����X�?             @       t       u                   @m@r�q��?             @       ������������������������       �                     @        v       w                 433�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        {       �                   `f@���.�d�?Z            �a@       |       }                   �h@�wY;��?X             a@        ������������������������       �        )            �P@        ~       �                    @L@�θV�?/            @Q@              �                   p`@�}�+r��?             C@       �       �       
             �?XB���?             =@       �       �                    �?h�����?             <@        �       �                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        �       �                   �`@�����H�?             "@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `@�חF�P�?             ?@       �       �                   @_@�q�q�?             8@       �       �                    �?��2(&�?             6@        ������������������������       �                      @        �       �                    �?R���Q�?             4@       �       �                    �?���!pc�?             &@       �       �                    �?�q�q�?             "@        �       �                   �]@z�G�z�?             @        ������������������������       �                     @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   n@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�Fǌ��?0            �S@        �       �                   �_@ 7���B�?             ;@        �       �                   @\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                     J@        �       �                    �?     ��?             0@        �       �                   �^@r�q��?             @        ������������������������       �                     @        �       �                   P`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �m@ s�n_Y�?              J@       �       �                    �?$��m��?             :@        �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@��.k���?             1@       �       �                    b@z�G�z�?             $@       �       �                    a@�����H�?             "@       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?$�q-�?             :@        �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@        �       �                   �[@�2�,��?(            �P@        ������������������������       �                     @        �       �                    �?�p����?#            �N@       �       �                    �?�LQ�1	�?             G@        �       �                     M@�����H�?             2@       ������������������������       �                     &@        �       �                    �?����X�?             @       �       �                    �N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ����?      �?             <@        ������������������������       �                      @        �       �                   �d@�z�G��?
             4@       �       �                   `c@z�G�z�?             .@       �       �                    �M@�z�G��?             $@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   `]@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   0d@������?             .@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  �"z?+�?���B`��?c��|��?s�3���?��T���?�K��T�?��Moz��?!Y�B�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?]t�E�?      �?      �?              �?      �?      �?              �?      �?                      �?ҏ~���?p�\��?����W�?�ѯz�@�?����k�?�5��P�?KKKKKK�?�������?      �?        ��,d!�?��Moz��?�������?�������?      �?              �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?      �?                      �?jv���*�?`�(tSR�?BE��f��?�{��ɣ?�D�)͋�?t�n���?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?      �?        �l�w6��?AL� &W�?              �?�E]t��?t�E]t�?      �?              �?      �?ffffff�?333333�?      �?      �?              �?�m۶m��?�$I�$I�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?      �?              �?              �?      �?      �?        t�E]t�?]t�E�?              �?      �?                      �?Cy�5��?^Cy�5�?^Cy�5�?(������?|���?>����?              �?      �?        �������?�������?              �?      �?        l(�����?(������?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        �B!��?��{���?h/�����?/�����?ZZZZZZ�?�������?      �?              �?      �?      �?      �?      �?      �?      �?                      �?              �?      �?        �������?�������?              �?      �?                      �?�Mozӛ�?�,d!Y�?�F��]�?-��>N��?��ٌ?I�dn�?r؃H{�?��6���?F]t�E�?]t�E�?�������?�������?      �?      �?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?6��9�?�]����?ZZZZZZ�?ZZZZZZ�?              �?�Q�g���?̵s���?(�����?�5��P�?�{a���?GX�i���?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?��RJ)��?�Zk����?�������?UUUUUU�?t�E]t�?��.���?              �?333333�?333333�?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?              �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�3���?1���M��?h/�����?	�%����?�������?�������?      �?                      �?              �?              �?      �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?;�;��?�;�;�?vb'vb'�?�N��N��?�q�q�?�q�q�?              �?      �?      �?              �?      �?        �?�������?�������?�������?�q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?              �?;�;��?�؉�؉�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?o�Wc"=�?"=P9���?              �?ާ�d��?C��6�S�?Nozӛ��?d!Y�B�?�q�q�?�q�q�?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?      �?      �?              �?ffffff�?333333�?�������?�������?ffffff�?333333�?      �?      �?      �?              �?      �?              �?      �?                      �?      �?        �������?333333�?      �?                      �?�?wwwwww�?�������?�������?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJB	VhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK�h��B�<         �                    �?4�5����?�           ��@               _                   �a@�.�0Q�?�            @w@                                  �?t���?�            �r@                                033�?     ��?             @@                                  �[@���Q��?             @        ������������������������       �                     �?               
       	             �?      �?             @               	                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                  �v@�����H�?             ;@                                 �U@$�q-�?             :@        ������������������������       �                     �?                                   @O@`2U0*��?             9@       ������������������������       �        	             0@                                  @L@�����H�?             "@                                  �?z�G�z�?             @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?               6                    �?l ��H|�?�            �p@               #                    �?��a�n`�?;            @W@                     
             �? ��WV�?#             J@        ������������������������       �                     5@                                  `_@`Jj��?             ?@        ������������������������       �                     ,@                                    �I@�t����?             1@        ������������������������       �                      @        !       "                   pe@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        $       +                    �?D^��#��?            �D@        %       &                    U@�G�z��?             4@        ������������������������       �                     �?        '       *                    �?D�n�3�?             3@       (       )                   �U@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ,       5                   �f@�G��l��?             5@       -       .                    �?j���� �?             1@        ������������������������       �                     @        /       4                    �?r�q��?             (@        0       3                   o@����X�?             @       1       2                    @I@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        7       X                    �?t���s��?o             f@       8       M                    @M@XI�~�?b            @c@       9       <                   @E@�d����?V            @a@        :       ;                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        =       F                    �?�\=lf�?T            �`@       >       ?       	             �?����}��?O            �_@        ������������������������       �        "             M@        @       E                   �a@@	tbA@�?-            @Q@        A       B                    �K@�IєX�?             1@       ������������������������       �        
             .@        C       D                 @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        !             J@        G       L                    �?؇���X�?             @       H       K       	             �?z�G�z�?             @        I       J                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        N       S                    �?     ��?             0@       O       P                   Pc@r�q��?	             (@       ������������������������       �                     "@        Q       R                   e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        T       U                    �M@      �?             @        ������������������������       �                      @        V       W                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Y       ^       	             �?\X��t�?             7@       Z       ]                 833�?X�<ݚ�?
             2@       [       \                 `ffֿz�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        `       g                    �L@��
P��?(            �Q@        a       d                    �D@�r����?             >@        b       c                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        e       f                   @g@$�q-�?             :@       ������������������������       �                     8@        ������������������������       �                      @        h       y                    �?      �?             D@       i       t                    �?�c�Α�?             =@       j       m                    �?������?             1@        k       l                    X@      �?             @        ������������������������       �                      @        ������������������������       �                      @        n       q                    �?8�Z$���?             *@       o       p                   �e@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        r       s                    c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       x       
             �?�q�q�?             (@       v       w                    �O@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        z       {                    �?"pc�
�?             &@        ������������������������       �                     �?        |                            N@ףp=
�?             $@        }       ~                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Y�*�?�            �v@        �       �                    �?��
ц��?'            @P@       �       �                 ����?��R[s�?            �A@        �       �                   pp@X�<ݚ�?             "@       �       �                   pe@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?8�Z$���?             :@       �       �       	             �?      �?             0@       �       �                    �?"pc�
�?             &@        ������������������������       �                      @        �       �                 ����?�<ݚ�?             "@       �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?z�G�z�?             $@        ������������������������       �                     @        �       �                     H@���Q��?             @        ������������������������       �                      @        �       �                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@�r����?             >@        �       �                    �?      �?             (@       �       �                    �?և���X�?             @        �       �                    b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@�X�<ݺ?             2@        �       �                    �I@r�q��?             @        �       �                   �k@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �? ��R��?�            �r@        �       �                    �?p�5�9��?N            �]@       �       �       
             �?�θ�?4            �S@       �       �                   �i@�S����?*            �L@        �       �                    �?     ��?             0@        �       �                    �?؇���X�?             @       �       �                    @M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   �\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?������?            �D@       �       �       	             �?��(\���?             D@       �       �                   �r@�X�<ݺ?             B@       �       �                    d@      �?             @@       ������������������������       �                     ;@        �       �                    �J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   pp@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �N@և���X�?
             5@       �       �                   �`@z�G�z�?             .@       �       �                   �q@�q�q�?             "@       �       �                    `@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?,���i�?            �D@       �       �                    �?��?^�k�?            �A@        �       �       
             �?��S�ۿ?
             .@       ������������������������       �                     *@        �       �                   `Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                   �n@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    a@�;Y�&��?v            @f@       �       �                   �[@�k.s�׌?\            �a@        �       �                   `[@���J��?"            �I@       ������������������������       �                     G@        �       �                   �`@z�G�z�?             @        ������������������������       �                     @        �       �                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        :            �V@        �       �                    �?���@��?            �B@        �       �                   b@      �?             $@        �       �                 ����?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �\@�����H�?             ;@        �       �                    �?      �?             @       �       �                   �n@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B0   Np	�?���Gw{�?P?���O�?`�X`�?G�#͑��?�q˸e�?      �?      �?333333�?�������?              �?      �?      �?      �?      �?              �?      �?              �?        �q�q�?�q�q�?;�;��?�؉�؉�?      �?        {�G�z�?���Q��?              �?�q�q�?�q�q�?�������?�������?              �?      �?      �?      �?                      �?              �?      �?        @�Ε$�?�6Ũ�o�?�c�1��?�s�9��?O��N���?;�;��?      �?        ���{��?�B!��?      �?        <<<<<<�?�?      �?        9��8���?�q�q�?      �?                      �?,Q��+�?�]�ڕ��?�������?�������?              �?l(�����?(������?;�;��?;�;��?              �?      �?                      �?1�0��?��y��y�?ZZZZZZ�?�������?      �?        UUUUUU�?�������?�$I�$I�?�m۶m��?�������?333333�?              �?      �?                      �?              �?      �?        3��Yb�?k��2�?5�wL��?V~B����?��\;0��?)�3J���?      �?      �?      �?                      �?"=P9���?g��1��?����~��?�@ �?      �?        �%~F��?ہ�v`��?�?�?      �?              �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?      �?              �?              �?      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?              �?      �?        !Y�B�?��Moz��?�q�q�?r�q��?�������?�������?              �?      �?                      �?      �?        PuPu�?_�_��?�������?�?      �?      �?      �?                      �?�؉�؉�?;�;��?      �?                      �?      �?      �?�{a���?5�rO#,�?�?xxxxxx�?      �?      �?              �?      �?        ;�;��?;�;��?F]t�E�?]t�E�?              �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?              �?      �?              �?        F]t�E�?/�袋.�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?����2��?A�ME��?�؉�؉�?�;�;�?X|�W|��?PuPu�?�q�q�?r�q��?UUUUUU�?�������?              �?      �?              �?        ;�;��?;�;��?      �?      �?/�袋.�?F]t�E�?      �?        9��8���?�q�q�?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�������?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?              �?�q�q�?��8��8�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?#�+��?��:\��?�O��O��?�����?�؉�؉�?ى�؉��?^Cy�5�?(������?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?������?�|����?333333�?�������?�q�q�?��8��8�?      �?      �?              �?�������?�������?              �?      �?              �?      �?              �?      �?              �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?              �?                      �?      �?        8��18�?�����?�A�A�?_�_��?�?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?��g<�?�0�9�a�?t�n��}?"����?�?______�?              �?�������?�������?              �?      �?      �?              �?      �?                      �?к����?L�Ϻ��?      �?      �?�������?UUUUUU�?              �?      �?                      �?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJMk/hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         h                    �?4�5����?�           ��@               ;                 ����?ٜSu��?�            �u@              6                    �?
�e4���?�             p@              	                   �O@�}�x�m�?�            �n@                                  `]@��
ц��?
             *@        ������������������������       �                     @                                   `Q@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        
       #                    �?`~A�P�?�             m@              "                   h@Pa�	�?y            �h@                     	             �?���p�T�?x            �h@                                   �?@-�_ .�?/            �R@                                 �t@F��}��?.            @R@                               ����? ��ʻ��?,             Q@                                  �G@���J��?"            �I@                                   �? �q�q�?             8@                                 @[@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     @        ������������������������       �                     ;@        ������������������������       �        
             1@                                  @`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                  �? �|ك�?I            �^@       ������������������������       �        F            @]@               !                    `@r�q��?             @                                   @L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        $       5                    �?4�2%ޑ�?            �A@       %       (                   �k@�LQ�1	�?             7@        &       '                   �a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        )       .                    �?�<ݚ�?             2@        *       +                     H@      �?             @        ������������������������       �                     �?        ,       -                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        /       0                 ����?؇���X�?             ,@        ������������������������       �                     "@        1       4                    �?���Q��?             @       2       3                    �H@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        7       8                   �_@      �?             (@        ������������������������       �                     @        9       :                    @M@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        <       _                    �?@�&b
}�?4            �U@       =       Z                   r@ޚ)�?*             R@       >       Y                   �o@�	j*D�?&            @P@       ?       P                 `ff@��}*_��?             K@       @       K                    �O@�G�z�?             D@       A       B                    ]@������?             A@        ������������������������       �                     "@        C       D                   h@`�Q��?             9@        ������������������������       �                     &@        E       F                     K@և���X�?             ,@        ������������������������       �                     @        G       H                    �?      �?              @       ������������������������       �                     @        I       J                     N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        L       M                   �\@r�q��?             @        ������������������������       �                     @        N       O                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Q       V                    �N@      �?             ,@       R       S                    
@      �?              @       ������������������������       �                     @        T       U                    �B@      �?             @        ������������������������       �                      @        ������������������������       �                      @        W       X                    �Q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        [       ^                 `ff�?����X�?             @        \       ]                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        `       e                    �?�r����?
             .@       a       d                    �J@$�q-�?             *@        b       c                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        f       g                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        i       �                    �?r=ά�{�?�            Px@        j       �                    �?
�K0��?[             a@       k       �                    �?������?D            �Y@       l       �                    �P@:~=�P�?6            @T@       m       �                    �?�(�Tw��?4            �S@       n       o                   �\@�iʫ{�?#            �J@        ������������������������       �                     @        p       {                   �_@�3Ea�$�?             G@        q       r                   @`@p�ݯ��?             3@        ������������������������       �                     @        s       x                    �?      �?             0@        t       u                    �?���Q��?             @        ������������������������       �                     �?        v       w                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                   �o@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        |       �                   l@�>����?             ;@        }       ~                   �d@"pc�
�?             &@       ������������������������       �                     @               �                    @C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        �       �                   �\@�q�����?             9@        ������������������������       �                     @        �       �                 ����?�eP*L��?             6@       �       �                    �?p�ݯ��?             3@       �       �                    b@ҳ�wY;�?	             1@       �       �                   @d@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �T@���7�?             6@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        �       �                     K@@�0�!��?             A@        �       �                   `\@      �?             (@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        �       �                   �e@�[|x��?�            �o@       �       �                   �a@ ��]��?�            `o@        ������������������������       �        %             M@        �       �                    �?��H���?{             h@       �       �                    �?M�D���?f            `c@        �       �                   �a@���|���?            �@@       �       �                   P`@�G��l��?             5@        �       �                    �?�q�q�?             (@        ������������������������       �                     �?        �       �                     J@���!pc�?             &@        �       �                    @H@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @O@�<ݚ�?             "@       �       �                   �a@      �?              @        �       �                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �H@�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �m@ @|���?P            �^@        �       �                   �m@ i���t�?#            �H@       �       �                   �X@=QcG��?"            �G@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   0m@`Ӹ����?             �F@       �       �                    �?��Y��]�?            �D@       �       �                   �\@���N8�?             5@        �       �                    �K@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �                     4@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   (q@��pBI�?-            @R@       �       �                    �?P���Q�?             D@       �       �                   0c@��?^�k�?            �A@       ������������������������       �                     @@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @z�G�z�?             @        ������������������������       �                      @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        �       �                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                     C@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP   Np	�?���Gw{�?s��\;0�?%~F���?���-iK�?�%mI[��?�z�����?�M!��?�؉�؉�?�;�;�?              �?۶m۶m�?�$I�$I�?      �?                      �?��x�w�?��� �?|���?|���?&���0�?J�f��?S�n0E�?к����?��Ǐ?�?����?�������?�?______�?�?�������?UUUUUU�?��y��y�?�a�a�?              �?      �?              �?              �?              �?        �������?333333�?      �?                      �?      �?        �_��e��?�h
���?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�A�A�?�������?d!Y�B�?Nozӛ��?�������?�������?      �?                      �?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?�������?333333�?      �?      �?      �?                      �?              �?              �?      �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        �C��:��?)^ ���?��8��8�?9��8���?;�;��?vb'vb'�?B{	�%��?_B{	�%�?�������?�������?�?xxxxxx�?              �?{�G�z�?��(\���?              �?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?      �?      �?                      �?�������?UUUUUU�?      �?                      �?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�?�؉�؉�?;�;��?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?0�;�O�?4=�,�?p�h�?n�?ȭ�;�H�?��;�o��?���O ��?�<ݚ�?��E���?�o��o��?� � �?
�[���?�琚`��?      �?        ����7��?��,d!�?^Cy�5�?Cy�5��?              �?      �?      �?�������?333333�?      �?              �?      �?      �?                      �?]t�E�?F]t�E�?      �?                      �?�Kh/��?h/�����?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?      �?        ���Q��?�p=
ף�?              �?t�E]t�?]t�E�?^Cy�5�?Cy�5��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?                      �?              �?F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?ZZZZZZ�?      �?      �?              �?      �?                      �?EQEQ�?]�u]�u�?ōOv�`�?G6q��?              �?�ҡ�3�?��+����?a�qa�?=���?F]t�E�?]t�E]�?1�0��?��y��y�?UUUUUU�?UUUUUU�?      �?        t�E]t�?F]t�E�?333333�?�������?              �?      �?                      �?9��8���?�q�q�?      �?      �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�}�K�`�?"XG��)�?����X�?/�����?AL� &W�?x6�;��?      �?      �?              �?      �?        l�l��??�>��?������?8��18�?�a�a�?��y��y�?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?      �?      �?      �?                      �?      �?        ����?���Ǐ�?�������?ffffff�?�A�A�?_�_��?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJH�_VhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKɅ�h��B@2         z                    �?�����?�           ��@              9                    �?h�T��v�?�            Px@                                  �a@0�n�"��?J             _@                                 �X@�����D�?(            @P@                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     @                                `ff@@�r-��?%            �M@       	                          �e@���5��?$            �L@       
                          �s@ �Cc}�?#             L@                                  �?�C��2(�?"            �K@                                  �`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                  @^@ "��u�?             I@                                   �?      �?             8@                                   �P@      �?              @                               ����?����X�?             @                                  `]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        ������������������������       �                     :@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �?L
�q��?"            �M@        ������������������������       �                     @                                    @B@���|���?            �K@        ������������������������       �                     @        !       8                    �?θ	j*�?             J@       "       +                    �?�\�u��?            �I@        #       $                   �]@ҳ�wY;�?             1@        ������������������������       �                     @        %       &                    �?��
ц��?             *@        ������������������������       �                      @        '       *                   `c@�eP*L��?             &@       (       )                   �k@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ,       7                    @J@�t����?             A@       -       0                    �E@���Q��?             9@        .       /       
             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        1       4                   Pd@���Q��?
             .@       2       3                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        5       6                   `g@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        :       o                    �?���s���?�            �p@       ;       d                    �?����?�            �j@       <       c                    �?H��2�?w            @g@       =       b                   �b@      �?S             `@       >       _                   �b@@4և���?I             \@       ?       R                    \@�IєX�?D            �Y@        @       O                    @�t����?             A@       A       F                    �?     ��?             @@        B       E                   �X@      �?              @        C       D                   @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        G       H                   �Y@�8��8��?             8@        ������������������������       �                     *@        I       J                   �k@"pc�
�?             &@       ������������������������       �                     @        K       L                   �Z@      �?             @        ������������������������       �                     �?        M       N                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        P       Q                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       V                    �?г�wY;�?/             Q@        T       U                     H@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �        
             ,@        W       X                    q@�O4R���?$            �J@       ������������������������       �                     B@        Y       Z                 `ff�?�IєX�?             1@       ������������������������       �                     *@        [       \                   @_@      �?             @        ������������������������       �                     �?        ]       ^                   `a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        `       a                 033�?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             0@        ������������������������       �        $             M@        e       f                    �?$�q-�?             :@        ������������������������       �                     @        g       h                    S@ףp=
�?             4@        ������������������������       �                     �?        i       j                    �?�}�+r��?             3@        ������������������������       �                     $@        k       l                   @a@�����H�?             "@       ������������������������       �                     @        m       n                    U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        p       s                    �J@^�!~X�?$            �J@        q       r                   `a@ҳ�wY;�?	             1@       ������������������������       �                     &@        ������������������������       �                     @        t       y                    �?������?             B@        u       v                   pc@$�q-�?
             *@       ������������������������       �                     &@        w       x                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        {       �                    �?0)RH'�?�            �u@       |       �                   h@4�ԗj�?�            �m@       }       �                    I@���+�ǲ?�            �m@        ~       �       	             �?և���X�?             @              �                   �a@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @O@0<�q �?�            �l@       �       �                   �?��wڝ�?~            @k@       ������������������������       �        g             f@        �       �                 033�?���N8�?             E@        �       �                    �?؇���X�?             ,@       �       �                    @L@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        �       �                   @t@���|���?             &@       �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����? ���]��?E            �Z@       �       �                    �?��ga�=�?.            �P@        �       �                    s@��S�ۿ?
             .@       ������������������������       �                     &@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �D@R�}e�.�?$             J@        �       �                    �?z�G�z�?             @       �       �                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @E@��[�p�?             �G@        �       �                    �?���!pc�?             &@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �      �?             @        ������������������������       �                     �?        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0d@�X�<ݺ?             B@       ������������������������       �                     :@        �       �                    �?z�G�z�?	             $@        ������������������������       �                     @        �       �                   �q@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�(�Tw��?            �C@        �       �                   �u@      �?
             0@       �       �                    �?�q�q�?	             .@        ������������������������       �                      @        �       �                    �?�θ�?             *@        �       �                     M@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   `c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @`@��<b���?             7@        ������������������������       �                     &@        �       �                   @b@�q�q�?             (@        ������������������������       �                     @        �       �                   ht@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  `�P47�?Њ�erd�?�"`�?�G7��g�?SJ)��R�?�Zk����?z�z��?z�z��?      �?      �?              �?      �?        ��c+���?'u_�?��Gp�?�}��?۶m۶m�?%I�$I��?F]t�E�?]t�E�?�������?333333�?      �?                      �?���Q��?�G�z�?      �?      �?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?                      �?              �?      �?              �?              �?        ��V'�?�pR���?      �?        ]t�E]�?F]t�E�?              �?�؉�؉�?�N��N��?�������?�?�������?�������?      �?        �;�;�?�؉�؉�?      �?        ]t�E�?t�E]t�?      �?      �?      �?                      �?      �?        �������?�������?333333�?�������?�������?�������?              �?      �?        �������?333333�?r�q��?�q�q�?      �?                      �?UUUUUU�?�������?      �?                      �?      �?                      �?q��;2l�?�a��y��?�V�9�&�?��`��}�?X`��?�~�駟�?      �?      �?�$I�$I�?n۶m۶�?�?�?�?<<<<<<�?      �?      �?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?F]t�E�?/�袋.�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�?�?�?�������?      �?                      �?�x+�R�?:�&oe�?              �?�?�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?              �?              �?;�;��?�؉�؉�?              �?�������?�������?      �?        (�����?�5��P�?              �?�q�q�?�q�q�?              �?      �?      �?      �?                      �?�	�[���?�}�	��?�������?�������?              �?      �?        �q�q�?�q�q�?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?              �?��k��?F��Q�g�?{CO��d�?M�[��?A�Iݗ��?��c+���?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?[9�\)�?����fԚ?N��ش�?�,�M�ɂ?      �?        ��y��y�?�a�a�?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?                      �?              �?      �?        ]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?                      �?��>���?Dj��V��?��[���?�1���?�������?�?      �?              �?      �?              �?      �?        'vb'vb�?�;�;�?�������?�������?      �?      �?      �?                      �?              �?�
br1�?m�w6�;�?t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ��8��8�?�q�q�?      �?        �������?�������?      �?        �m۶m��?�$I�$I�?      �?                      �?� � �?�o��o��?      �?      �?UUUUUU�?UUUUUU�?      �?        �؉�؉�?ى�؉��?�$I�$I�?�m۶m��?              �?      �?        UUUUUU�?�������?              �?      �?              �?        ��Moz��?��,d!�?              �?�������?�������?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	NhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK酔h��B@:         `                   �`@T8���?�           ��@               /                    �?�θ�?�            �u@               
                    �?��؇>��?V            @`@               	                    �?���B���?             :@                                   �?      �?             $@                                 �\@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             0@                                   �?�E��
��?G             Z@                                  �?�^����?'            �M@                                   �?�q�q�?             @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  �h@ �h�7W�?#            �J@       ������������������������       �                     @@                                   �?؇���X�?             5@                                  �E@ףp=
�?             4@        ������������������������       �                     �?                                `ff�?�}�+r��?             3@                                   �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?               *                    �?�<ݚ�?             �F@              )                    �?������?            �B@              "                    �E@ >�֕�?            �A@                !                   �\@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        #       $                    �?      �?             @@       ������������������������       �                     6@        %       &                 @33�?ףp=
�?             $@       ������������������������       �                      @        '       (                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        +       .                    �?      �?              @        ,       -                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        0       =                    �?�!/�'�?�            �k@        1       4                   �]@���?            �D@       2       3                    `Q@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        5       :                   �_@�\��N��?             3@        6       9                    �?z�G�z�?             $@       7       8                   @a@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ;       <                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        >       G                    �?`Ӹ����?j            �f@        ?       F                    �?��Y��]�?.            �T@        @       A                   �]@�q�q�?             @        ������������������������       �                      @        B       E                    �?      �?             @       C       D                   0o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        *             S@        H       Q                    `@��<D�m�?<            �X@        I       J                   �Y@PN��T'�?             ;@        ������������������������       �                     $@        K       L                   �[@������?             1@        ������������������������       �                     @        M       P                    \@@4և���?	             ,@        N       O                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        R       S                   `a@�J�T�?+            �Q@        ������������������������       �                     :@        T       _                    �?`Ӹ����?            �F@       U       V                    �?@-�_ .�?            �B@        ������������������������       �                     &@        W       ^                    `@$�q-�?             :@       X       Y                    @K@`2U0*��?             9@       ������������������������       �        	             *@        Z       ]                    �?�8��8��?             (@        [       \                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        a       �                    �?R�7�o�?�            �w@       b       �                    �?��a�2��?�             k@        c       �                   0e@     ��?,             P@       d       e                 ����?���3L�?%             K@        ������������������������       �                     @        f                           �P@r�qG�?              H@       g       z                    @f.i��n�?            �F@       h       k                    \@���"͏�?            �B@        i       j                    �M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        l       u                    @K@     ��?             @@       m       n                   e@ףp=
�?             4@        ������������������������       �                     �?        o       p                 ����?�}�+r��?             3@       ������������������������       �                     &@        q       r                    �?      �?              @        ������������������������       �                     �?        s       t                   @_@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        v       y                    �M@�q�q�?
             (@       w       x                   Pl@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        {       ~                   �`@      �?              @        |       }                   �\@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �B@z�G�z�?             $@        ������������������������       �                     �?        �       �                   �k@�����H�?             "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   h@�}�+r��?e             c@       �       �                   �?`2U0*��?d            �b@       �       �                    �O@P����?P            �]@       �       �                    �? �O�H�?K            �[@        ������������������������       �                     :@        �       �                   @[@`��>�ϗ?7            @U@        ������������������������       �                     �?        ������������������������       �        6             U@        �       �                   pa@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @@        ������������������������       �                     $@        �       �                   pa@"pc�
�?             6@        ������������������������       �                     @        �       �                   @b@      �?	             0@        ������������������������       �                      @        �       �       	             �?؇���X�?             ,@        �       �                   �k@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?����d�?b            �d@       �       �                    �?>�b���?M            @`@       �       �                    �?�%o��?(            �P@        �       �                   �a@���Q��?             4@       �       �                   y@��S���?	             .@       �       �                    �?�n_Y�K�?             *@        �       �                    �L@؇���X�?             @        ������������������������       �                      @        �       �                 033@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   0c@�7����?            �G@       �       �                    �?z�G�z�?             D@        �       �                   �m@�n_Y�K�?             *@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�����H�?             ;@        �       �                    b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?ףp=
�?             4@       ������������������������       �                     .@        �       �                    U@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   pd@����X�?             @        ������������������������       �                     @        �       �                    \@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@���N8�?%            �O@        �       �                   �i@$�q-�?             :@        ������������������������       �                     (@        �       �                     M@؇���X�?	             ,@       ������������������������       �                     &@        �       �                    �O@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Hq@^H���+�?            �B@       �       �                   �j@�θ�?             :@        �       �                    �C@      �?              @        ������������������������       �                     �?        �       �                   �d@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    \@�X�<ݺ?             2@        �       �                    �L@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        �       �                     K@���|���?             &@        ������������������������       �                     @        �       �                    @M@z�G�z�?             @        ������������������������       �                      @        �       �                   �s@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�L���?            �B@       ������������������������       �                     >@        �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                 833�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  6n����?�� ���?�؉�؉�?ى�؉��??�?��?�~�~�?��؉���?ى�؉��?      �?      �?�$I�$I�?�m۶m��?              �?      �?              �?              �?        ��؉���?;�;��?W'u_�?u_[4�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        "5�x+��?��sHM0�?              �?�$I�$I�?۶m۶m�?�������?�������?      �?        (�����?�5��P�?UUUUUU�?�������?              �?      �?                      �?      �?        9��8���?�q�q�?��g�`��?к����?��+��+�?�A�A�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?���ٴ?=�d=�d�?8��18�?28��1�?F]t�E�?�.�袋�?              �?      �?        �5��P�?y�5���?�������?�������?�m۶m��?�$I�$I�?              �?      �?              �?        �q�q�?�q�q�?      �?                      �?l�l��??�>��?������?8��18�?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?և���X�?��S�r
�?h/�����?&���^B�?              �?�?xxxxxx�?      �?        �$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?��V؜?(�K=�?              �?l�l��??�>��?к����?S�n0E�?              �?;�;��?�؉�؉�?{�G�z�?���Q��?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?��b����?�&:�Bd�?��8��8�?�q�q�?     ��?      �?�%���^�?&���^B�?              �?�������?�������?�`�`�?�>�>��?v�)�Y7�?*�Y7�"�?�������?333333�?              �?      �?              �?      �?�������?�������?              �?�5��P�?(�����?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?              �?              �?�������?�������?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?              �?�5��P�?(�����?���Q��?{�G�z�?�V'u�?'u_[�?c��2��?5'��Ps�?      �?        �������?�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?        /�袋.�?F]t�E�?      �?              �?      �?              �?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?              �?      �?              �?                      �?S&���?�l��4�?�����?~�~��?\�՘H�?���[��?�������?333333�?�?�������?;�;��?ى�؉��?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?G}g����?]AL� &�?�������?�������?ى�؉��?;�;��?      �?                      �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?              �?�������?333333�?      �?                      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �a�a�?��y��y�?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        L�Ϻ��?�g�`�|�?ى�؉��?�؉�؉�?      �?      �?      �?        �$I�$I�?�m۶m��?      �?                      �?��8��8�?�q�q�?�������?�������?      �?                      �?      �?        F]t�E�?]t�E]�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        L�Ϻ��?}���g�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���%hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�7         f                    �?�����?�           ��@              %                    �?�D�e�?�?�            pw@                                  �?4�ԗj�?�            �m@                                ���@�Z��L��?-            �Q@                                  �?���7�?+            �P@                                 `c@����˵�?(            �M@       ������������������������       �        #            �J@               	                     J@      �?             @        ������������������������       �                     �?        
                           �?���Q��?             @                                  �?      �?             @                                 �e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?�Ń��̧?e             e@                                   �?�q�q�?             @                                  @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               $                    �? �Jj�G�?b            �d@                                  @L@ � ���?\            �c@                                 @[@ 
�V�?O            �`@                      
             �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        J            �^@                !                   Hp@�8��8��?             8@       ������������������������       �        
             1@        "       #                     M@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        &       5                    �?��.k���?Y             a@        '       ,                    �?z�G�z�?            �A@       (       )                   �]@��s����?             5@        ������������������������       �                     $@        *       +                   �T@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        -       0                    �?d}h���?
             ,@        .       /                   �W@      �?             @        ������������������������       �                      @        ������������������������       �                      @        1       4                   @\@ףp=
�?             $@        2       3                   �[@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       S                    �?�7�yHx�?A            @Y@       7       L                 ����?�J�T�?/            �Q@       8       9                 `ffֿP̏����?'            �L@        ������������������������       �                      @        :       ;                    �?�rF���?%            �K@        ������������������������       �                     $@        <       I                    �?������?            �F@       =       B                    @F@<ݚ)�?             B@        >       ?                   `]@և���X�?	             ,@        ������������������������       �                     @        @       A                   pf@      �?              @       ������������������������       �                     @        ������������������������       �                      @        C       D                    �L@��2(&�?             6@       ������������������������       �                     1@        E       F                    �?���Q��?             @        ������������������������       �                     �?        G       H                   �b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        J       K                   @Y@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        M       R                   0a@X�Cc�?             ,@       N       Q                    �?"pc�
�?             &@       O       P                   �[@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        T       e                    �?�z�G��?             >@       U       V                   `_@��.k���?             1@        ������������������������       �                     @        W       X                    �?      �?	             (@        ������������������������       �                     @        Y       Z                    ]@�q�q�?             "@        ������������������������       �                     �?        [       b                    �?      �?              @       \       ]                   `b@z�G�z�?             @        ������������������������       �                      @        ^       _                    �?�q�q�?             @        ������������������������       �                     �?        `       a                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        c       d                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        g       �                    �?���҅�?�            pv@        h       s                    �F@�lwd2V�?P            �`@        i       r                   �a@�q�q�?             8@       j       q                    �?���N8�?             5@       k       l                    �?�IєX�?             1@        ������������������������       �                     @        m       n                   �o@�C��2(�?             &@       ������������������������       �                      @        o       p       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        t       �                   p`@�G�.o�?A            @[@        u       |                    �?�LQ�1	�?             G@        v       {                    �?r�q��?             @       w       z       	             �?      �?             @       x       y                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        }       ~                 ����?��Q���?             D@        ������������������������       �                     (@               �       
             �?��>4և�?             <@        �       �                    @��
ц��?             *@       �       �                    �L@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@�q�q�?             .@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �                    `@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��s����?'            �O@       �       �                    @�I�w�"�?             C@       �       �                   0k@�z�G��?             >@        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                   @a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��s����?             5@        �       �                 `ff�?և���X�?             @       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                      @        �       �                    �?H%u��?             9@       �       �                    �?      �?             (@        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@       ������������������������       �                     @        �       �                     M@      �?             @        ������������������������       �                     �?        �       �                    �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?4��Q���?�            @l@       �       �                   0f@nS޸��?i             f@        ������������������������       �                     ?@        �       �                    �?��W��?V            @b@        �       �                    @O@      �?             0@       �       �                    �?�n_Y�K�?             *@       �       �                    �?X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   @_@      �?              @        ������������������������       �                      @        �       �                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?8�Z$���?K            @`@        �       �                    �?��<D�m�?            �H@        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                   �Z@�(\����?             D@        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �B@        �       �                   @h@.�	F�9�?/            @T@        �       �                   �g@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                    ]@>A�F<�?,             S@        �       �                    �?��S���?             .@       �       �                    @I@�eP*L��?             &@        �       �                   0o@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �K@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    @M@Xny��?%            �N@       �       �                    @K@ �q�q�?             H@       ������������������������       �                    �@@        �       �                   �m@�r����?             .@        �       �                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        �       �                   @b@�n_Y�K�?	             *@       �       �                   �Z@�����H�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        (            �H@        �t�b�`     h�h)h,K ��h.��R�(KK�KK��hi�B�  ������?�v
��,�?�E�����?y�&1��?{CO��d�?M�[��?���.�d�?��Vؼ?�.�袋�?F]t�E�?W'u_�?��/���?      �?              �?      �?      �?        �������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?                      �?��<��<�?�a�a�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        k߰�k�?��)A��?ɞ��td�?�&��jq�?������?g��1�~?]t�E�?F]t�E�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �m۶m��?�$I�$I�?              �?      �?              �?        �?�������?�������?�������?�a�a�?z��y���?              �?F]t�E�?]t�E]�?      �?                      �?۶m۶m�?I�$I�$�?      �?      �?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?#
L:5�?��g����?H���@��?p�z2~��??���#�?��Gp�?              �?yJ���?�־a��?      �?        wwwwww�?�?��8��8�?�8��8��?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?��.���?t�E]t�?      �?        �������?333333�?              �?      �?      �?      �?                      �?�q�q�?�q�q�?              �?      �?        �m۶m��?%I�$I��?F]t�E�?/�袋.�?�������?�������?      �?                      �?      �?              �?        333333�?ffffff�?�������?�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?mR�ګ�?�+E	��?�RKE,�?�VwZ�i�?UUUUUU�?UUUUUU�?�a�a�?��y��y�?�?�?      �?        ]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��p�?z|���?d!Y�B�?Nozӛ��?�������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?333333�?              �?I�$I�$�?۶m۶m�?�؉�؉�?�;�;�?۶m۶m�?�$I�$I�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �a�a�?z��y���?�5��P�?����k�?333333�?ffffff�?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �a�a�?z��y���?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?              �?              �?���Q��?)\���(�?      �?      �?      �?        F]t�E�?/�袋.�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?x�!���?����	�?�^o�?�?G($��?              �?Ĉ#F��?ϝ;w���?      �?      �?;�;��?ى�؉��?�q�q�?r�q��?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?;�;��?;�;��?և���X�?��S�r
�?�q�q�?9��8���?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?~X�<��?�����H�?333333�?�������?              �?      �?        Cy�5��?������?�������?�?]t�E�?t�E]t�?�������?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?        �}�K�`�?C��6�S�?UUUUUU�?�������?              �?�?�������?      �?      �?      �?                      �?              �?ى�؉��?;�;��?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJs-hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKӅ�h��B�4         �       
             �?>�����?�           ��@                     	             �?�f���?b           (�@              @                    �?�^��&
�?�            0y@                                   �?*�~�9��?b            �a@                                   �?ܷ��?��?             =@        ������������������������       �                     @                                  `c@ȵHPS!�?             :@                               ����?�nkK�?	             7@       	                           @N@ףp=
�?             $@        
                           �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�\��N��?V            �\@                                   x@ �Cc}�?             <@       ������������������������       �                     9@        ������������������������       �                     @               -                    �?֦�r��?B            �U@                                  �D@��0u���?,             N@                                  �a@X�<ݚ�?	             "@        ������������������������       �                      @                                   �B@����X�?             @                                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               $                    P@������?#            �I@                #                    �?����X�?             @        !       "                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        %       &                    d@fP*L��?             F@       ������������������������       �                     :@        '       (                    @I@b�2�tk�?             2@        ������������������������       �                     @        )       *                    _@�q�q�?             (@        ������������������������       �                     @        +       ,                   f@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        .       /                   �^@�	j*D�?             :@        ������������������������       �                     @        0       ?                    b@�ՙ/�?             5@       1       2                    �?������?             1@        ������������������������       �                     �?        3       >                 `ff�?      �?             0@       4       =                     M@z�G�z�?             .@       5       6                    `@�q�q�?             "@        ������������������������       �                     �?        7       8                   �d@      �?              @       ������������������������       �                     @        9       :                    a@�q�q�?             @        ������������������������       �                     �?        ;       <                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        A       P                    �?H�8���?�            @p@        B       E                 ����?d}h���?             <@        C       D                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        F       G                 833�?r�q��?             8@        ������������������������       �                     @        H       O                   b@���y4F�?             3@        I       J                    ]@      �?              @        ������������������������       �                     �?        K       N                     L@և���X�?             @       L       M                    Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        Q       T                   @Z@�NI���?�             m@        R       S                   �Y@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        U       `                    �?F��}��?�            `k@        V       W                   �k@��`qM|�?0            �T@       ������������������������       �                     G@        X       Y                    �?������?            �B@        ������������������������       �                     &@        Z       ]                   pm@8�Z$���?             :@        [       \                   @_@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ^       _                   �e@�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        a       b                    �?�IєX�?R             a@        ������������������������       �                     @        c       j                    @K@���}��?Q            �`@        d       i                    @G@P����?&            �M@        e       f                    �?�}�+r��?             3@       ������������������������       �        
             1@        g       h                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     D@        k       ~                   �a@�����?+            �R@       l       o                    �K@:�&���?            �C@        m       n                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        p       }                 `ff @4?,R��?             B@       q       r                   �i@z�G�z�?             9@       ������������������������       �                     *@        s       v                    `@�q�q�?             (@        t       u                 tff�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        w       |                   `b@�q�q�?             "@       x       {                    �?؇���X�?             @        y       z                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                    �A@        �       �                 pff�?�+I�9��?f            @f@       �       �                 ����? �\���?Y            �c@       �       �                   p@�J�T�?Q            �a@       ������������������������       �        2             X@        �       �                    �?���}<S�?             G@       �       �                    �?t��ճC�?             F@       �       �                   `p@��Y��]�?            �D@        �       �                 @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     C@        �       �                   �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �\@      �?             0@        ������������������������       �                     @        �       �                   Pt@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                   Pr@���Q��?             4@       �       �                    �?�t����?             1@        ������������������������       �                     @        �       �                   d@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�X���x�?`             c@       �       �                 033�?xP�Fֺ�?7            @V@       �       �                    �O@ ��Ou��?1            �S@       �       �                    �?xL��N�?.            �R@       �       �                   �b@ ��ʻ��?+             Q@        ������������������������       �                     A@        �       �                 @33�?г�wY;�?             A@       �       �                   �n@`2U0*��?             9@        �       �                   �\@�����H�?             "@        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        ������������������������       �                     "@        �       �                 033�?�q�q�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    п      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �I@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �F@     ��?)             P@        ������������������������       �                     @        �       �                   P`@0B��D�?$            �M@        �       �                    �N@     ��?             @@       �       �                   Pk@�<ݚ�?             ;@       ������������������������       �                     .@        �       �                   �?      �?             (@        ������������������������       �                     @        �       �                    �?؇���X�?             @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?PN��T'�?             ;@        �       �                    �Q@���!pc�?	             &@       ������������������������       �                     @        �       �                    k@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �`@      �?
             0@       ������������������������       �                     $@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  ���� �?u(���o�?�������?"�%��?�c��)
�?"N�	���?�L[����?fI9 2�?��=���?a���{�?      �?        ��N��N�?�؉�؉�?�Mozӛ�?d!Y�B�?�������?�������?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�5��P�?y�5���?۶m۶m�?%I�$I��?              �?      �?        ��/���?���/��?�������?""""""�?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?xxxxxx�?�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?颋.���?]t�E]�?      �?        �8��8��?9��8���?      �?        �������?�������?      �?              �?      �?              �?      �?        ;�;��?vb'vb'�?              �?�a�a�?�<��<��?�?xxxxxx�?              �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?              �?        �J��J��?�Vj�Vj�?۶m۶m�?I�$I�$�?      �?      �?              �?      �?        UUUUUU�?�������?              �?(������?6��P^C�?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?              �?���=��?��FX��?�؉�؉�?ى�؉��?              �?      �?        ����?��Ǐ?�?��k���?�@	o4u�?              �?к����?��g�`��?              �?;�;��?;�;��?۶m۶m�?�$I�$I�?              �?      �?        (�����?�5��P�?              �?      �?        �?�?              �?���̮?4�τ?�?'u_[�?�V'u�?(�����?�5��P�?              �?      �?      �?      �?                      �?              �?v�)�Y7�?�Ϻ���?�o��o��?�A�A�?UUUUUU�?UUUUUU�?      �?                      �?r�q��?�8��8��?�������?�������?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?              �?�3��g�?�as�ü?���7a�?�3���?(�K=�?��V؜?      �?        ӛ���7�?d!Y�B�?�E]t��?t�E]t�?8��18�?������?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?      �?      �?              �?�؉�؉�?;�;��?      �?                      �?�������?333333�?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        �)�)�?W�W��?�.p��?�я~���?.��-���?�i�i�?>�S��?L�Ϻ��?�������?�?      �?        �?�?���Q��?{�G�z�?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?t�E]t�?      �?                      �?      �?      �?      �?        ��}ylE�?�A�I��?      �?      �?�q�q�?9��8���?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?        h/�����?&���^B�?t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�E^hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKͅ�h��B@3         |                    �?F���?��?�           ��@              E                    �?V�-Vz�?           �z@              2                    �?���_���?�            �p@                                   �?V�K/��?2            �S@                                  �?Fx$(�?             I@                                   �?������?	             1@              
                 ����?�r����?             .@               	                   `b@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                      	             �?"pc�
�?            �@@                                  �?HP�s��?             9@                                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?���7�?             6@                                   @N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@                                   @C@      �?              @        ������������������������       �                     @                                   �?z�G�z�?             @                                   �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @               +                   �o@����"�?             =@              "                    `@      �?             4@                !                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #       *                    �?@�0�!��?             1@       $       )                    @d}h���?
             ,@       %       (                   �?�8��8��?             (@        &       '                    @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ,       -                    �L@�q�q�?             "@        ������������������������       �                      @        .       1                   xq@؇���X�?             @        /       0                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        3       D                    �?�q�q��?y             h@       4       5                    �?�ȨF=�?q            `f@        ������������������������       �        $            �K@        6       7                    @G@�&/�E�?M             _@        ������������������������       �                    �K@        8       C                   Pg@�θV�?/            @Q@       9       :                   n@t�e�í�?.            �P@       ������������������������       �                    �C@        ;       >                   @[@�>4և��?             <@        <       =                   @c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ?       @                   �?���}<S�?             7@       ������������������������       �                     3@        A       B                   xp@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        F       _                    �?��Q���?b             d@        G       H                 ����?�5U��K�?0            �T@        ������������������������       �                    �A@        I       ^                   {@r�q��?             H@       J       Q                 ����?��0{9�?            �G@        K       L                    @I@�q�q�?             @        ������������������������       �                     �?        M       N                    �?z�G�z�?             @        ������������������������       �                     �?        O       P                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        R       [                   pc@��p\�?            �D@       S       Z                    `@�7��?            �C@        T       Y                   �^@�r����?             .@       U       X                    �?@4և���?             ,@       V       W                    @Q@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        \       ]                   pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        `       y                    �?"+q��?2            @S@       a       n                    �?�d�����?)            �L@       b       g                 ����?�r����?             �F@       c       f                    X@��?^�k�?            �A@        d       e                 @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @@        h       m                    �?      �?             $@       i       j                   0l@����X�?             @        ������������������������       �                     @        k       l                   �_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        o       x                    `P@      �?	             (@       p       w                   �f@"pc�
�?             &@       q       v                 @33�?ףp=
�?             $@       r       u                    d@�����H�?             "@        s       t                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        z       {                   `\@z�G�z�?	             4@       ������������������������       �                     0@        ������������������������       �                     @        }       �                   �a@R��jf��?�            �r@       ~       �       	             �?��[�8��?�            �i@              �                   Pf@�YTV��?z            �g@        �       �                   �`@������?*             R@       ������������������������       �        $            �N@        �       �                   �`@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �J@t�I��n�?P            @]@        �       �       
             �?H�z�G�?             D@       �       �                   i@^������?            �A@        �       �                    �B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?������?             >@       �       �                    �?d}h���?             <@       �       �                   `j@�㙢�c�?             7@        �       �                   �i@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�����H�?             2@       �       �                    �?      �?             0@       �       �                   �\@��S�ۿ?             .@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?j(���?3            @S@        �       �                 ����?��
ц��?             :@        �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 hff�?�����?             3@        ������������������������       �                      @        �       �                    �M@ҳ�wY;�?             1@       �       �                   `W@d}h���?	             ,@        ������������������������       �                     �?        �       �                    �?8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @        �       �                   �a@���J��?!            �I@       ������������������������       �                     F@        �       �                   �j@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?	             .@        �       �                   j@r�q��?             @        �       �                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �       
             �?Pa�	�?>            �X@       �       �                   �`@����?�?9            �V@       �       �                    �R@(;L]n�?'             N@       �       �                 033�?P����?&            �M@        �       �                    �?���7�?             6@        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                    �B@        ������������������������       �                     �?        ������������������������       �                     >@        �       �                    �M@�����H�?             "@        ������������������������       �                     @        �       �                   ``@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ,�U�)�?js���?�R��}�?�Z�c(�?�ެ'�6�?@�La�$�?�Z܄��?�ґ=�?R���Q�?ףp=
��?xxxxxx�?�?�������?�?9��8���?�q�q�?      �?                      �?      �?                      �?F]t�E�?/�袋.�?{�G�z�?q=
ףp�?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        	�=����?�i��F�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?ZZZZZZ�?�������?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?UUUUU��?�������?�R"x���?���}��?      �?        2�c�1�?�s�9�?      �?        ̵s���?�Q�g���?�1����?�rv��?      �?        �$I�$I�?�m۶m��?�������?333333�?              �?      �?        ӛ���7�?d!Y�B�?      �?              �?      �?              �?      �?                      �?      �?        �������?333333�?��k���?���h��?              �?UUUUUU�?�������?L� &W�?m�w6�;�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?      �?                      �?��+Q��?�]�ڕ��?�A�A�?��[��[�?�?�������?�$I�$I�?n۶m۶�?;�;��?�؉�؉�?              �?      �?                      �?      �?                      �?      �?      �?      �?                      �?      �?        �wL��?�g�'��?Cy�5��?y�5���?�������?�?_�_��?�A�A�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?              �?              �?      �?F]t�E�?/�袋.�?�������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?              �?        �������?�������?              �?      �?        pu�8���?�"�1K	�?�������?�?lp����?壓�N>�?�q�q�?�q�q�?              �?F]t�E�?/�袋.�?      �?                      �?���?�s?�s?�?333333�?ffffff�?_�_��?uPuP�?�������?�������?              �?      �?        �?wwwwww�?۶m۶m�?I�$I�$�?d!Y�B�?�7��Mo�?�������?333333�?              �?      �?        �q�q�?�q�q�?      �?      �?�?�������?      �?      �?              �?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?�������?333333�?              �?      �?              �?              �?        ��cj`��?�g�'��?�;�;�?�؉�؉�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?Q^Cy��?^Cy�5�?      �?        �������?�������?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?      �?                      �?              �?�?______�?              �?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        |���?|���?l�l��?��I��I�?�?�������?'u_[�?�V'u�?F]t�E�?�.�袋�?      �?                      �?              �?      �?                      �?�q�q�?�q�q�?              �?�������?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�&UhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK�h��B�<         6                    �F@"�\�&U�?�           ��@               %                    �?�I�w�"�?^             c@                                  �?��Õty�?F             ]@        ������������������������       �                     @                                    �?��X��?C             \@                                  �?�X�<ݺ??             [@                                  �?`�(c�?8            �X@        ������������������������       �                     0@        	                           _@Ћ����?-            �T@        
                           ^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �?�Fǌ��?+            �S@        ������������������������       �        
             3@                                   l@ �.�?Ƞ?!             N@                     
             �?�nkK�?             7@                                  @D@$�q-�?             *@                                  �C@؇���X�?             @       ������������������������       �                     @                                  pf@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                    �B@                                  �_@�z�G��?             $@                                  �?      �?             @                                   C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        !       "                    �?      �?             @        ������������������������       �                     �?        #       $       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        &       5       
             �?*O���?             B@       '       0                   �^@�������?             >@        (       -                    �?և���X�?
             ,@        )       ,                    �E@����X�?             @       *       +                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        .       /                     E@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        1       2       	             �?      �?             0@       ������������������������       �        	             ,@        3       4                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        7       �                    �?b���L��?l           0�@        8       g                    �?�^`���?�            �l@       9       >                    �?W@e��?k            �c@        :       =                    a@�eP*L��?             &@       ;       <                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ?       Z                   �d@��ӄ���?c            @b@       @       W                    �?|�9ǣ�?Q            �]@       A       J                    �?p���h�?J            @[@        B       I       	             �?�(\����?             D@       C       D                   �b@�nkK�?             7@       ������������������������       �                     4@        E       H                    �?�q�q�?             @       F       G                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        K       L                   �?�θV�?/            @Q@       ������������������������       �        !            �G@        M       P                   Pi@�X����?             6@        N       O                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        Q       R                   `a@      �?             (@        ������������������������       �                     @        S       V       	             �?؇���X�?             @       T       U                    a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        X       Y                    V@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        [       b                    �?����X�?             <@        \       a                    �?      �?              @       ]       ^                   �^@���Q��?             @        ������������������������       �                      @        _       `       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        c       f                   0k@R���Q�?             4@        d       e                    j@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        h       �                    �?�E����?0             R@       i       j                    �?Hث3���?            �C@        ������������������������       �                     "@        k       n                    �?d��0u��?             >@        l       m                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        o       ~                    �?�q�q�?             ;@       p       }                   �p@      �?             0@       q       x                    �?�q�q�?             (@        r       w                   �b@����X�?             @       s       t                   �_@      �?             @        ������������������������       �                     �?        u       v                   @m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        y       |                 `ff�?���Q��?             @        z       {                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               �                   pj@�eP*L��?             &@       �       �                    V@      �?              @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �R@�C��2(�?            �@@       �       �                     K@      �?             @@        �       �       
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ;@        ������������������������       �                     �?        �       �                    �?pס���?�            v@        �       �                   �c@ ��/K��?F            �Z@       �       �                 ����? ��~���?;            �V@        �       �                   �b@�?�|�?            �B@       ������������������������       �                     B@        ������������������������       �                     �?        �       �                    �Q@�T`�[k�?&            �J@       �       �                    �?Jm_!'1�?"            �H@        �       �                 ����?�eP*L��?             &@        ������������������������       �                     @        �       �                   �p@      �?              @       �       �                    @N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�˹�m��?             C@       �       �                   0b@�X�<ݺ?             B@       ������������������������       �                     8@        �       �                    �?r�q��?
             (@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �       
             �?���Q��?             @        ������������������������       �                     �?        �       �                   Pb@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	             �?      �?             0@       �       �                    �N@�eP*L��?             &@       �       �                   @n@؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �J@$�q-�?�            �n@        �       �                    @J@؇���X�?"             L@       �       �                    �?Hm_!'1�?            �H@        �       �                    �I@և���X�?             @       �       �                    �H@z�G�z�?             @       �       �                    b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @G@�Ń��̧?             E@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     B@        �       �                   �\@և���X�?             @        ������������������������       �                     @        �       �                   �l@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ����? �r�ɻ?i            �g@        �       �       
             �?�?�<��?"            @P@       �       �                    �?�X�<ݺ?             K@       �       �                     P@     ��?             @@       �       �                   �`@��2(&�?             6@        �       �                    _@�q�q�?             @        ������������������������       �                     @        �       �                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@      �?
             0@        �       �                    �?�����H�?             "@        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        	             6@        �       �                     L@�eP*L��?             &@        ������������������������       �                      @        �       �                   `l@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    r@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�Ń��̧?G            �_@        �       �                    �?$�q-�?             :@       ������������������������       �                     7@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    c@ �ׁsF�?8             Y@       ������������������������       �        4            �W@        �       �                    @N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  ��j��`�?:�J;�O�?����k�?�5��P�?�FX�i�?��=���?              �?۶m۶m�?%I�$I��?��8��8�?�q�q�?��)x9�?և���X�?      �?        ԮD�J��?��+Q��?UUUUUU�?UUUUUU�?              �?      �?        1���M��?�3���?      �?        wwwwww�?�?�Mozӛ�?d!Y�B�?�؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?              �?              �?        ffffff�?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?�������?�������?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        �:*���?����?Ψ5����?e����f�?�9A��?A����?t�E]t�?]t�E�?۶m۶m�?�$I�$I�?              �?      �?                      �?_�z����?�
*T��?Jݗ�V�?�A�Iݷ?l�O����?�,�M�ɲ?333333�?�������?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?        ̵s���?�Q�g���?      �?        �E]t��?]t�E]�?�������?�������?      �?                      �?      �?      �?      �?        �$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?333333�?�$I�$I�?۶m۶m�?      �?                      �?      �?        �q�q�?r�q��?�i�i�?��-��-�?      �?        wwwwww�?DDDDDD�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?]t�E�?t�E]t�?      �?      �?�������?333333�?              �?      �?                      �?      �?        F]t�E�?]t�E�?      �?      �?�������?333333�?      �?                      �?              �?      �?        ��|u�?=,�P1�?�}�	��?�`��}�?�'}�'}�?�`�`�?к����?*�Y7�"�?              �?      �?        "5�x+��?���!5��?������?����X�?t�E]t�?]t�E�?      �?              �?      �?UUUUUU�?�������?      �?                      �?      �?        ^Cy�5�?��P^Cy�?�q�q�?��8��8�?              �?UUUUUU�?�������?�q�q�?9��8���?              �?�������?333333�?      �?              �?      �?      �?                      �?              �?      �?      �?              �?      �?              �?      �?      �?              �?      �?      �?                      �?      �?      �?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?              �?        ;�;��?�؉�؉�?�$I�$I�?۶m۶m�?9/���?Y�Cc�?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �a�a�?��<��<�?UUUUUU�?�������?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?              �?      �?                      �?o��2�|�?�ќ5(�? �����?�����?�q�q�?��8��8�?      �?      �?t�E]t�?��.���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?              �?]t�E�?t�E]t�?              �?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?                      �?�a�a�?��<��<�?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?{�G�z�?�G�z��?              �?�������?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�uhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKυ�h��B�3         j                    �?R������?�           ��@              M                    �?�+�o�?�?�            �w@                                 @E@(��+�?�            s@               	                    �?l��[B��?             =@                      	             �?�n_Y�K�?             *@                                  �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        
                           �?     ��?             0@                                  �?ףp=
�?             $@                      	             �?�q�q�?             @                                  �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?��ś��?�            @q@                                   �?      �?             (@                                  �?�eP*L��?             &@                                  �J@r�q��?             @                      
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               J                   h@(�B'�?�            �p@               +                    \@��{$h�?�            0p@        !       &                 tff�?H�V�e��?             A@       "       #                   @c@ �Cc}�?             <@        ������������������������       �                     ,@        $       %                   �c@d}h���?
             ,@        ������������������������       �                     @        ������������������������       �        	             &@        '       *                   �[@�q�q�?             @       (       )                     M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ,       5                    @L@���
���?�             l@       -       .                    �?�B:�g�?k            �e@       ������������������������       �        Y            @b@        /       0                 433�?h�����?             <@       ������������������������       �                     6@        1       4                   �`@r�q��?             @        2       3                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       G                    s@L紂P�?!            �I@       7       >                    b@�:�^���?            �F@       8       =                   �_@г�wY;�?             A@        9       :                   �o@r�q��?             @       ������������������������       �                     @        ;       <       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        ?       F                    �?���!pc�?             &@       @       A                    �?�����H�?             "@        ������������������������       �                     @        B       C                    m@z�G�z�?             @        ������������������������       �                     @        D       E                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        H       I                 ����?      �?             @        ������������������������       �                     @        ������������������������       �                     @        K       L                   pn@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        N       O                    �?h/��y��?2            @S@        ������������������������       �                     @        P       c                   �o@z��R[�?,            �Q@       Q       b       	             �?�5��
J�?             G@       R       _                   �b@�<ݚ�?            �F@       S       ^                 ��� @�KM�]�?             C@       T       ]                    m@�㙢�c�?             7@       U       \                    �?��2(&�?             6@       V       [                    c@�θ�?	             *@       W       X                    �?r�q��?             (@        ������������������������       �                     @        Y       Z                 `ff�?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        
             .@        `       a                 033�?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        d       e                    �?�8��8��?             8@       ������������������������       �        	             0@        f       i                   a@      �?              @        g       h                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        k       �       	             �?��!pc�?�             v@       l       �                    �?�LQ�1	�?�             t@        m       t                    _@�	j*D�?6            �S@        n       q                   �a@�û��|�?             7@        o       p                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        r       s                 ����?@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        u       �                   @q@"pc�
�?'            �K@       v       w                    \@�q��/��?#            �H@        ������������������������       �                     "@        x       �                   0n@R���Q�?             D@       y       �                   0m@�n`���?             ?@       z                           �?�����H�?             ;@       {       ~                 pff�?���N8�?             5@        |       }                     R@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             (@        �       �                   �]@�q�q�?             @        ������������������������       �                     �?        �       �                   �c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   Pm@      �?             @       �       �                    @P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    @L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �e@�٠n�}�?�            �n@       �       �                   ``@������?�            `n@        �       �                    �O@�?�'�@�?L            �\@       �       �                    �?4��?�?G             Z@        �       �                   �r@�n_Y�K�?             *@       �       �                    �?X�<ݚ�?             "@       �       �                     I@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?0�>���??            �V@       �       �                    @�g<a�?5            @S@       �       �                    �?�k~X��?1             R@        ������������������������       �                     (@        �       �                 033�? �.�?Ƞ?)             N@       ������������������������       �                    �@@        �       �                   `_@ 7���B�?             ;@       ������������������������       �        	             0@        �       �                   @`@�C��2(�?             &@        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �H@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �]@d}h���?
             ,@        �       �                   �]@���Q��?             @        ������������������������       �                     �?        �       �                   �X@      �?             @        ������������������������       �                     �?        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�����H�?             "@        �       �                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @]@      �?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@ g�yB�?M             `@        �       �                   @b@ ��WV�?             J@       ������������������������       �                     G@        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        �       �                   �c@z�G�z�?             @        ������������������������       �                     @        �       �                 @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        /            @S@        ������������������������       �                     �?        �       �                   �b@���Q��?             >@       �       �                    @L@�	j*D�?             :@       �       �                    W@�����H�?
             2@        ������������������������       �                      @        ������������������������       �        	             0@        �       �                   �k@      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b��(     h�h)h,K ��h.��R�(KK�KK��hi�B�  ��*��?5��j���?_�%���?B��U@�?q�����?;ڼOq��?GX�i���?���=��?ى�؉��?;�;��?�������?�������?      �?                      �?      �?              �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?R�g���?s��\;0�?      �?      �?t�E]t�?]t�E�?�������?UUUUUU�?      �?      �?              �?      �?              �?        �������?�������?      �?                      �?              �?��&�l��?m��&�l�?Y�	R�%�?q�a�
��?iiiiii�?ZZZZZZ�?%I�$I��?۶m۶m�?      �?        I�$I�$�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?2Tv����?߼�xV4�?��f���?Ȥx�L�w?      �?        �m۶m��?�$I�$I�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?}�'}�'�?l�l��?�?�?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        F]t�E�?t�E]t�?�q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?      �?                      �?              �?      �?      �?              �?      �?        �������?�������?      �?                      �?V~B����?���15��?      �?        X|�W|��?���?�Mozӛ�?�,d!Y�?�q�q�?9��8���?(�����?�k(���?d!Y�B�?�7��Mo�?t�E]t�?��.���?�؉�؉�?ى�؉��?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?      �?              �?                      �?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?              �?      �?                      �?�E]t��?�.�袋�?Y�B��?��Moz��?;�;��?vb'vb'�?8��Moz�?��,d!�?�q�q�?�q�q�?      �?                      �?n۶m۶�?�$I�$I�?              �?      �?        F]t�E�?/�袋.�?և���X�?/����?              �?333333�?333333�?�c�1��?�9�s��?�q�q�?�q�q�?�a�a�?��y��y�?�q�q�?�q�q�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?      �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �u�y��?Pq����?�:���?�������?y�5���?������?ى�؉��?�N��N��?ى�؉��?;�;��?r�q��?�q�q�?      �?      �?              �?      �?              �?                      �?�!�!�?��=��=�?�cj`?���8+�?�q�q�?�8��8��?              �?�?wwwwww�?              �?h/�����?	�%����?              �?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?�������?�������?      �?                      �?۶m۶m�?I�$I�$�?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        ����?�����?;�;��?O��N���?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?      �?                      �?              �?      �?        333333�?�������?vb'vb'�?;�;��?�q�q�?�q�q�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�G5GhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�7         �       	             �?<���m�?�           ��@              u                   �b@��E��V�?s           �@              "                    �?��oh���?           `{@                                  0d@�fSO��?A            �X@                                  �e@�+$�jP�?             ;@                                  �Q@8�Z$���?             :@              
                 ������8��8��?             8@               	                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                      @        ������������������������       �                     �?                                   �?��ӭ�a�?/             R@                                  �?�q�q�?'             N@                                  �?@-�_ .�?            �B@       ������������������������       �                    �@@                                  �b@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                hff�?��<b���?             7@        ������������������������       �                     "@                                    L@X�Cc�?             ,@        ������������������������       �                     @                                   �?X�<ݚ�?             "@        ������������������������       �                     @                                  �\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @               !                 ����?�8��8��?             (@                                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        #       H                    �?>��i3�?�            0u@        $       5                    �?�Pf����?;            �W@        %       2                    �?�^�����?            �E@       &       )                    �?@�0�!��?             A@        '       (                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        *       /                    `P@��� ��?             ?@       +       .                   @E@`2U0*��?             9@        ,       -                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        0       1                   `a@      �?             @        ������������������������       �                     @        ������������������������       �                     @        3       4                   �R@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        6       E                   �r@D>�Q�?"             J@       7       D                    �?��E�B��?            �G@        8       C                   pm@      �?             0@       9       >                   �_@���Q��?             .@       :       =                   �]@؇���X�?             @        ;       <                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ?       B                    b@      �?              @       @       A                   @`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ?@        F       G                   �^@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        I       ^                    �?`R�
�?�            �n@        J       [                    �?�חF�P�?             ?@       K       Z                    �?ȵHPS!�?             :@       L       Y                   b@@�0�!��?
             1@       M       P                    �?�z�G��?             $@        N       O                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Q       R                    �?      �?              @        ������������������������       �                     �?        S       T                   @`@����X�?             @        ������������������������       �                     �?        U       X                   @m@r�q��?             @        V       W                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        \       ]                     M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        _       h                   `_@�J�T�?�            �j@       `       a                    �?`��(�?U            �`@        ������������������������       �        "            �M@        b       c                    �?P�Lt�<�?3             S@        ������������������������       �                     4@        d       e                   �k@h�����?%             L@       ������������������������       �                     A@        f       g                    �?�C��2(�?             6@        ������������������������       �                      @        ������������������������       �                     4@        i       n                   `@�7��?0            �S@        j       m                    �?�θ�?             *@       k       l                    @L@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        o       p                    �? ����?(            @P@       ������������������������       �        !             K@        q       r                    �?�C��2(�?             &@        ������������������������       �                     @        s       t                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        v       {                   �Q@���w��?_            �a@        w       x                 033@$�q-�?             *@       ������������������������       �                     &@        y       z                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       �                    �?     x�?X             `@       }       �                    �?�0���?:            �T@       ~       �                    �?�q��/��?              G@              �                   Pd@ >�֕�?            �A@        �       �                    �?      �?
             0@       �       �                 @33�?@4և���?             ,@        �       �                    �?�����H�?             "@       �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    �N@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        �       �                    �?���!pc�?             &@       ������������������������       �                     @        �       �                 833@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                   Pd@��+��?            �B@        �       �                   �c@�E��ӭ�?             2@        ������������������������       �                     @        �       �                     M@�r����?
             .@        �       �                    �?      �?             @       �       �                   �m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?�d�����?             3@        ������������������������       �                     @        �       �                    �H@�q�q�?             .@       �       �                    @F@z�G�z�?             $@       �       �                   pf@����X�?             @       �       �                   �e@r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @K@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�ݏ^���?            �F@       �       �                    �?��Zy�?            �C@        �       �                    �?      �?	             0@       �       �                   �g@�C��2(�?             &@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �t@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?\X��t�?             7@       �       �                   �_@��S���?             .@       �       �                   �c@      �?              @        ������������������������       �                     �?        �       �                   �e@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �q@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �H@      �?              @        ������������������������       �                     @        �       �                    �N@      �?             @       �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? Ņ殲�?a            `c@       �       �                    �? qP��B�?Q             `@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                   e@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �P@ ��7��?N            �^@        �       �                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        K            @]@        �       �                   �o@      �?             :@        �       �                   �^@z�G�z�?             .@        ������������������������       �                     @        ������������������������       �                     (@        �       �                     J@�C��2(�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ���>��?�,@��"�?���,��??;��i�?����?ȏ?~��?�v�ļ�?w�ļ�!�?B{	�%��?/�����?;�;��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        ��8��8�?�8��8��?UUUUUU�?UUUUUU�?S�n0E�?к����?      �?              �?      �?      �?                      �?��Moz��?��,d!�?              �?�m۶m��?%I�$I��?              �?r�q��?�q�q�?      �?        �������?�������?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?�.�	��?�{���G�?a�+F�?�-q����?�5eMYS�?֔5eMY�?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?              �?      �?        �{����?�B!��?���Q��?{�G�z�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?�q�q�?9��8���?      �?                      �?vb'vb'�?b'vb'v�?AL� &W�?�l�w6��?      �?      �?�������?333333�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?333333�?�������?      �?                      �?�����??�%C���?��RJ)��?�Zk����?�؉�؉�?��N��N�?�������?ZZZZZZ�?333333�?ffffff�?      �?      �?              �?      �?              �?      �?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?              �?�������?333333�?              �?      �?        ��V؜?(�K=�?t��:W�?j�����?              �?(�����?���k(�?              �?�$I�$I�?�m۶m��?              �?F]t�E�?]t�E�?      �?                      �?�A�A�?��[��[�?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?                      �? �����? �����?              �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?���=��?i^���S�?;�;��?�؉�؉�?              �?      �?      �?              �?      �?             ��?      �?o4u~�!�?"�%��?�B����?��Mozӻ?��+��+�?�A�A�?      �?      �?n۶m۶�?�$I�$I�?�q�q�?�q�q�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?              �?        F]t�E�?t�E]t�?      �?        �������?333333�?      �?                      �?�S�n�?*�Y7�"�?r�q��?�q�q�?      �?        �?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?Cy�5��?y�5���?      �?        UUUUUU�?UUUUUU�?�������?�������?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        ��I��I�?�[�[�?� � �?\��[���?      �?      �?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        �������?333333�?              �?      �?        ��Moz��?!Y�B�?�������?�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?��%�_��?mЦm�?��}A�?�}A_З?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        ��:ڼ�?;ڼOqɀ?�������?�������?              �?      �?              �?              �?      �?�������?�������?              �?      �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJO�#hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         p                 ����?8}�ý�?�           ��@              !                   `@LМ_���?�             x@                                   �?�kwY���??            @Z@                                   �?H.�!���?             I@        ������������������������       �                      @                                ����?     ��?             H@                                  �?���H��?             E@                                  �?$�q-�?            �C@       	       
                    `Q@�g�y��?             ?@       ������������������������       �                     >@        ������������������������       �                     �?                                    P@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �?�q�q�?             @                                 `X@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                   @K@,�+�C�?             �K@        ������������������������       �                     :@                                  �k@\-��p�?             =@        ������������������������       �        
             ,@                                    �?������?
             .@                                  �?���Q��?             $@                                   L@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        "       9                    �?@���e��?�            �q@        #       $                    �?r٣����?'            �P@        ������������������������       �                      @        %       4                    n@     ��?%             P@       &       3       	             �?P����?             C@       '       .                    �?r�q��?             >@       (       )                 ����?PN��T'�?             ;@       ������������������������       �                     5@        *       +                    �?�q�q�?             @        ������������������������       �                      @        ,       -                   0m@      �?             @        ������������������������       �                      @        ������������������������       �                      @        /       2                    �?�q�q�?             @       0       1                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        5       6                 833�? ��WV�?             :@       ������������������������       �                     8@        7       8       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        :       _                    �?�ʈD��?�            �j@       ;       @                    P@����!p�?o             f@        <       ?                    �?      �?             @        =       >                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        A       X                   �?!�;��?k            �e@       B       W       	             �?Kb8�į?b            �c@       C       T                   �b@xdQ�m��?2            @T@       D       Q                    �M@�7��?0            �S@       E       L                    �?��pBI�?,            @R@       F       G                    @G@�\=lf�?)            �P@       ������������������������       �                    �B@        H       K                   �c@(;L]n�?             >@       I       J                   �b@@4և���?             ,@       ������������������������       �        
             *@        ������������������������       �                     �?        ������������������������       �                     0@        M       P                   �d@r�q��?             @       N       O       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        R       S                    �P@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        U       V                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        0            �R@        Y       Z                    �?      �?	             0@        ������������������������       �                     @        [       ^                 pff�?r�q��?             (@        \       ]                   @a@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        `       c                   �j@��Sݭg�?            �C@        a       b       	             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        d       g                    �?6YE�t�?            �@@        e       f                   �r@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        h       k                    q@��s����?             5@       i       j                    \@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        l       m                   �^@      �?             @        ������������������������       �                     �?        n       o                    �H@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        q       �                    �?t���-��?�            �u@       r       �                 `ff @v�|����?�            0r@       s       �                    �?�rF���?�            �k@       t       �                   pa@z�G�z�?�            @j@       u       v                   �[@L`EU�P�?e            �b@        ������������������������       �                     �I@        w       �                    �P@B�1V���?E            @X@       x       }                    �? 	��p�??            �U@        y       z                    �?և���X�?             @        ������������������������       �                     @        {       |                     F@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                 ����?x�G�z�?9             T@               �                    �?�KM�]�?             3@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                    �?��v$���?,            �N@        �       �       
             �?(;L]n�?             >@       �       �                   �T@P���Q�?             4@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     $@        ������������������������       �                     ?@        �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Xr@V{q֛w�?&             O@       �       �                    �?䯦s#�?             �J@       �       �                   �`@��
ц��?            �C@       �       �                    �?���Q��?             9@       �       �                    �?�eP*L��?             6@       �       �       
             �?d}h���?             ,@        ������������������������       �                     @        �       �                     J@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                     J@      �?              @        �       �                    @E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	             �?d}h���?             ,@       �       �                    d@8�Z$���?             *@       ������������������������       �                     "@        �       �                   �X@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?؇���X�?             ,@       ������������������������       �                     "@        �       �                   �`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                 ����?���Q��?             $@        ������������������������       �                     @        �       �                   0n@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @L@ ��PUp�?,            �Q@        �       �                   c@�C��2(�?             &@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        &             N@        �       �       
             �?F�����?$            �L@       �       �                    @K@��S���?            �F@        �       �                 ����?@�0�!��?             1@       ������������������������       �                     $@        �       �                     E@և���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 033�?      �?             <@       �       �                    �?      �?
             0@        �       �                   �k@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                 033@      �?             (@       �       �                     P@؇���X�?             @        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    U@r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  a[ӿc�?PR Np�?�'b6��?j�;����?Z�5Z�5�?S.�R.��?�(\����?)\���(�?              �?      �?      �?�0�0�?��y��y�?�؉�؉�?;�;��?��{���?�B!��?      �?                      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?��)A��?�}��7��?              �?�{a���?a����?              �?�?wwwwww�?�������?333333�?      �?      �?      �?                      �?      �?                      �?�(�I�?�\����?|���?>���>�?      �?              �?      �?Q^Cy��?�P^Cy�?UUUUUU�?�������?h/�����?&���^B�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        ;�;��?O��N���?              �?      �?      �?      �?                      �?A_���?�}A_з?/�袋.�?]t�E�?      �?      �?      �?      �?      �?                      �?              �?�)kʚ��?6eMYS֤?�o��o��?�i�i�?�5?,R�?X�<ݚ�?��[��[�?�A�A�?���Ǐ�?����?"=P9���?g��1��?      �?        �������?�?n۶m۶�?�$I�$I�?      �?                      �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        �|˷|��?�i�i�?UUUUUU�?�������?              �?      �?        '�l��&�?e�M6�d�?UUUUUU�?UUUUUU�?      �?                      �?z��y���?�a�a�?�������?�?              �?      �?              �?      �?      �?        �������?333333�?      �?                      �?��֡�l�?�L�Ȥ�?��ǿ���?[P���?�־a��?yJ���?�������?�������?#�u�)�?L�Ϻ��?              �?��4l7��?���$2�?�{a���?������?۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?        333333�?�������?(�����?�k(���?UUUUUU�?UUUUUU�?      �?                      �?              �?;ڼOqɐ?.�u�y�?�?�������?�������?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?�������?�������?      �?              �?      �?      �?                      �?�{����?B!��?�V�9�&�?�����?�؉�؉�?�;�;�?333333�?�������?t�E]t�?]t�E�?I�$I�$�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?      �?        ۶m۶m�?I�$I�$�?;�;��?;�;��?              �?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?�������?333333�?      �?                      �?9��8���?�q�q�?      �?                      �?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?��V،?��ۥ���?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?              �?u�YLg�?�YLg1�?�������?�?ZZZZZZ�?�������?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?              �?      �?              �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?�������?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��^hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�=         �                    �?�����?�           ��@                                  �?`�X�?           �{@                      	             �?d/
k�?D             [@                                 `c@�� =[�?,             Q@                                  �?��a�n`�?(             O@                                  �? �h�7W�?#            �J@       ������������������������       �                     E@               	                   �R@���!pc�?
             &@        ������������������������       �                      @        
                           �?�����H�?	             "@       ������������������������       �                     @                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  @V@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @                      
             �?r�q��?             @                                ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     D@               �       	             �?Ԑ ̽�?�            �t@              l                    �?a��t��?�            @m@              -                   �]@      �?r             f@               $                    �?�4�����?             ?@               #                    f@      �?
             $@              "                    �?      �?              @              !                     I@���Q��?             @                                  `^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        %       &                    �?���N8�?             5@       ������������������������       �                     (@        '       ,                    �K@X�<ݚ�?             "@       (       +                   �[@r�q��?             @       )       *                    e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        .       _                 033�?8^s]e�?Y             b@       /       L                   (p@z�G�z�?K             ^@       0       C                    �?H�g�}N�?7            �V@       1       @                   �f@���(-�?+            @R@       2       ;                 833�?�J�T�?)            �Q@       3       :                    �? ����?%            @P@       4       5                   d@���J��?            �I@       ������������������������       �                    �@@        6       9       
             �?�X�<ݺ?
             2@        7       8                    �I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     ,@        <       ?       
             �?r�q��?             @       =       >                    a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        A       B                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       K                   0m@      �?             2@       E       F                    �K@���Q��?             .@        ������������������������       �                     @        G       J                   �a@      �?              @       H       I                    �O@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        M       V                    �G@�f7�z�?             =@        N       U                   �c@؇���X�?             ,@        O       T                   �x@����X�?             @       P       Q                    �?r�q��?             @        ������������������������       �                     @        R       S                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        W       ^                   q@�q�q�?             .@        X       [                    �?      �?              @        Y       Z                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        \       ]                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        `       a                    �?�J�4�?             9@        ������������������������       �                     "@        b       k                   pm@      �?             0@       c       h                    �?X�<ݚ�?             "@       d       g                    �?�q�q�?             @       e       f                   �h@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        i       j                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        m       z       
             �?^l��[B�?(             M@       n       q                    �?��S�ۿ?            �F@        o       p                     Q@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        r       w                    �?�IєX�?             A@       s       t                    �? ��WV�?             :@       ������������������������       �                     7@        u       v                   `\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        x       y                   `@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        {       �                    �?�θ�?	             *@       |                        @33�?      �?              @        }       ~                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    _@���Q��?             @        ������������������������       �                      @        �       �                    �P@�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `X@`{��T��?9            @Y@        ������������������������       �                     @        �       �                    @�)���Y�?8            �X@       �       �                   �g@�8��8N�?7             X@       �       �                    �?��	,UP�?5             W@       �       �                   �?(;L]n�?4            �V@       ������������������������       �        *            �P@        �       �                    @L@      �?
             8@       ������������������������       �                     2@        �       �                    �L@      �?             @        ������������������������       �                      @        �       �                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �h@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?v�|����?�            0r@       �       �                    �?�����	�?�            �o@        �       �                    �?�eP*L��?             6@       �       �                   �a@$�q-�?	             *@       ������������������������       �                     $@        �       �                   `b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?h�{��`�?�             m@        �       �                   �s@����X�?             <@       �       �                   `c@r�q��?             8@       �       �                    �?������?             .@       �       �                   @m@8�Z$���?
             *@        �       �                    �G@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?���(��?�            �i@       �       �                   (q@h�[F���?a            `b@       �       �                 ����?Ԫ2��?K            �\@        �       �                   �i@      �?             D@        ������������������������       �                     2@        �       �                   �d@�eP*L��?             6@       �       �                    �?���Q��?             4@        �       �                 ����?r�q��?             @        �       �                   `m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   0j@      �?             ,@        ������������������������       �                     @        �       �                     J@���|���?             &@       �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�L���?2            �R@        �       �                   @`@z�G�z�?             .@        ������������������������       �                     @        �       �                   �`@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @G@����˵�?&            �M@        �       �                   �Z@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                    @M@@�E�x�?!            �H@       ������������������������       �                     ?@        �       �                   Pa@�X�<ݺ?             2@       ������������������������       �                     $@        �       �                    a@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �@@        �       �                    �?XB���?&             M@       �       �                    _@������?            �D@       ������������������������       �                     6@        �       �                    �?�KM�]�?             3@       �       �                    �H@�r����?	             .@        �       �                    �?���Q��?             @       �       �                    �      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     1@        �       �                    �?*O���?             B@       �       �                    �?�������?             >@       �       �                    �?p�ݯ��?             3@       �       �                    c@����X�?             ,@       �       �                    ]@r�q��?             (@        ������������������������       �                     @        �       �                   �r@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   `@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  `�P47�?Њ�erd�?N[R�?�cI��[�?�Kh/���?/�����?�������?�������?�s�9��?�c�1Ƹ?��sHM0�?"5�x+��?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        �yO�0@�?�a/��?!� ��?��[��[�?      �?      �?��RJ)��?���Zk��?      �?      �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ��y��y�?�a�a�?              �?r�q��?�q�q�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?|a���?	�=����?�������?�������?|��{���?���?��իW��?�P�B�
�?(�K=�?��V؜? �����? �����?______�?�?      �?        ��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?              �?      �?�������?333333�?              �?      �?      �?      �?      �?              �?      �?              �?              �?        O#,�4��?a���{�?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?              �?{�G�z�?�z�G��?              �?      �?      �?�q�q�?r�q��?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?��=���?�=�����?�?�������?F]t�E�?]t�E�?              �?      �?        �?�?;�;��?O��N���?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        ى�؉��?�؉�؉�?      �?      �?      �?      �?      �?                      �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?!w�l�2�?�F�tj�?              �?Dc}h��?������?�������?�������?d!Y�B�?��Mozӫ?�������?�?      �?              �?      �?      �?              �?      �?              �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?                      �?��ǿ���?[P���?�?{{{{{{�?]t�E�?t�E]t�?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        >����?�n�	�m�?�$I�$I�?�m۶m��?UUUUUU�?�������?�?wwwwww�?;�;��?;�;��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        z�gaz�?1=ӳ0�?���+ݻ?!͎Z��?p�}��?$���>��?      �?      �?              �?]t�E�?t�E]t�?�������?333333�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?        F]t�E�?]t�E]�?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        L�Ϻ��?}���g�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?��/���?W'u_�?�������?�������?      �?                      �?9/���?և���X�?              �?�q�q�?��8��8�?              �?      �?      �?              �?      �?                      �?�{a���?GX�i���?������?p>�cp�?              �?(�����?�k(���?�?�������?�������?333333�?      �?      �?              �?      �?                      �?              �?              �?              �?�q�q�?�q�q�?�������?�������?Cy�5��?^Cy�5�?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?      �?              �?        333333�?�������?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�	�^hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�Mh�h)h,K ��h.��R�(KM��h��B�@         �                    �?.��X~��?�           ��@                                  �?�����?           �y@                                   �?Υf���?(            �N@                      
             �?��a�n`�?             ?@               
                   �`@X�Cc�?	             ,@                                  �?      �?              @        ������������������������       �                      @               	                     G@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                ����?�t����?
             1@                                 �b@�<ݚ�?             "@                                 �m@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �J@z�G�z�?             >@                                  @[@���Q��?             $@        ������������������������       �                      @                                   �?      �?              @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@                W                    �?�mqA{��?�            �u@        !       B                   �b@�LQ�1	�?@             W@       "       A                 `ff�?�z�6�?)             O@       #       :                    �?r�qG�?             H@       $       )       
             �?�θ�?            �C@        %       (                   @j@���Q��?             .@        &       '                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        *       7                    �?      �?             8@       +       6                    �?�C��2(�?             6@       ,       3                   �`@ףp=
�?             4@       -       .                    �?�X�<ݺ?             2@        ������������������������       �                     @        /       2                     N@�C��2(�?             &@        0       1                     K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        4       5                    n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        8       9                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ;       >                    �?X�<ݚ�?             "@       <       =                    b@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ?       @       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        C       P                    @d��0u��?             >@       D       M                   Xq@���N8�?             5@       E       L                 ����?�t����?             1@       F       K                    �?"pc�
�?	             &@        G       J                    �?���Q��?             @       H       I                   e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        N       O                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        Q       R                 `ff@�q�q�?             "@        ������������������������       �                     @        S       V                    �?���Q��?             @       T       U                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        X       �                    `R@�?�            �o@       Y       p                    �?�X�<ݺ?�            �o@        Z       g                   ``@Xny��?+            �N@       [       \                    �?�}�+r��?             C@       ������������������������       �                     2@        ]       d                    �?ףp=
�?             4@       ^       _                 ����?�X�<ݺ?             2@        ������������������������       �                      @        `       a                   hq@ףp=
�?	             $@       ������������������������       �                      @        b       c                    @L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       f                   �h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        h       o                   pv@��<b���?             7@       i       n                   �i@"pc�
�?             6@       j       m                     M@���Q��?             $@        k       l                 ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     �?        q       |                    �?���q��?r            �g@        r       {                 ����?�Ń��̧?/             U@        s       t                   �i@ 	��p�?             =@       ������������������������       �        
             3@        u       z                   �`@z�G�z�?             $@        v       y                   `Z@      �?             @       w       x                   (q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �K@        }       ~                   �U@�f�¦ζ?C            �Z@        ������������������������       �                     �?               �                    `@�&=�w��?B            �Z@        �       �                   �_@��p\�?            �D@       �       �                    \@�}�+r��?             C@       �       �                    �?�C��2(�?             6@       �       �                    �I@"pc�
�?             &@       ������������������������       �                      @        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        
             0@        �       �                   �m@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @M@ ����?)            @P@       ������������������������       �                    �C@        �       �                    �? ��WV�?             :@       ������������������������       �        	             0@        �       �                    �M@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?��絹�?�            `t@       �       �                    �K@J�yE�?�            �o@       �       �                   @g@(.�`(�?m             e@       �       �       	             �?��`qM|�?l            �d@       �       �                   �[@��y� �?<            @W@        �       �                    �G@      �?             4@       �       �                    �C@      �?             $@        ������������������������       �                     @        �       �                 ���������X�?             @        ������������������������       �                     �?        �       �                    \@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?���(-�?/            @R@        ������������������������       �        
             0@        �       �                    �?�}�+r��?%            �L@       �       �                    @K@ 7���B�?"             K@       �       �                   �f@@�E�x�?            �H@       ������������������������       �                    �D@        �       �                    �?      �?              @        ������������������������       �                      @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        0            @R@        ������������������������       �                     @        �       �                 833�?8�$�>�?-            �U@       �       �                    �O@�{r٣��?"            �P@       �       �       	             �?`��}3��?            �J@       �       �                    �?F�����?            �F@       �       �       
             �?p9W��S�?             C@       �       �                    �?� �	��?             9@       �       �                    i@և���X�?             5@        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                   @b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             (@       �       �                    �?���!pc�?             &@        �       �                    �M@�q�q�?             @        ������������������������       �                     �?        �       �                   �i@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    ^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �^@$�q-�?             *@        �       �                    ]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?P���Q�?             4@       �       �                     N@��S�ۿ?             .@        �       �                   �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    U@R_u^|�?.            �Q@        �       �                     M@�q�q�?             8@       ������������������������       �        	             .@        �       �                    �?X�<ݚ�?             "@        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @a@      �?             @       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �                           �?�*/�8V�?             �G@       �       �                    �?�(�Tw��?            �C@       �       �                    @M@�>����?             ;@       ������������������������       �                     5@        �       �       
             �?�q�q�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?	             (@       �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                 ����?      �?             @        ������������������������       �                     �?        �       �                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KMKK��hi�B0  ��� ���?���o���?xxxxxx�?�������?.�u�y�?i�>�%C�?�c�1��?�s�9��?%I�$I��?�m۶m��?      �?      �?      �?        �������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?<<<<<<�?�?9��8���?�q�q�?      �?      �?      �?                      �?              �?      �?        �������?�������?333333�?�������?              �?      �?      �?      �?      �?              �?      �?        �������?UUUUUU�?      �?                      �?              �?)��п��?6��В�?d!Y�B�?Nozӛ��?�Zk����?J)��RJ�?UUUUUU�?UUUUUU�?�؉�؉�?ى�؉��?�������?333333�?      �?      �?      �?                      �?              �?      �?      �?F]t�E�?]t�E�?�������?�������?�q�q�?��8��8�?              �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�q�q�?r�q��?333333�?�������?              �?      �?              �?      �?      �?                      �?              �?DDDDDD�?wwwwww�?�a�a�?��y��y�?<<<<<<�?�?/�袋.�?F]t�E�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�������?�q�q�?��8��8�?�}�K�`�?C��6�S�?(�����?�5��P�?              �?�������?�������?�q�q�?��8��8�?              �?�������?�������?              �?      �?      �?      �?                      �?      �?      �?              �?      �?        ��Moz��?��,d!�?F]t�E�?/�袋.�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �]Ɣ�â?#�����?�a�a�?��<��<�?�{a���?������?              �?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?�Ե��?��4>2��?      �?        �x+�R�?tHM0���?��+Q��?�]�ڕ��?(�����?�5��P�?F]t�E�?]t�E�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?         �����? �����?              �?;�;��?O��N���?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?e@=S���?n�
�E�?�������?�������?��t����?8�Z$���?�@	o4u�?��k���??���O?�?X`��?      �?      �?      �?      �?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?      �?        ��իW��?�P�B�
�?      �?        �5��P�?(�����?	�%����?h/�����?և���X�?9/���?      �?              �?      �?      �?        �������?UUUUUU�?      �?                      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?6eMYS��?�5eMYS�?��|��?|���?�琚`��?M0��>��?�>�>��?؂-؂-�?�k(����?l(�����?�Q����?)\���(�?�$I�$I�?۶m۶m�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        �������?�������?      �?                      �?      �?              �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?�������?�������?�?      �?      �?              �?      �?              �?              �?        �@�6�?2~�ԓ��?�������?UUUUUU�?              �?r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?                      �?�٨�l��?AL� &W�?�o��o��?� � �?�Kh/��?h/�����?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJR��zhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         ~                    �?z��K���?�           ��@              a       
             �?�������?           �y@                                  �?H�` |�?�            pt@                                   �?���|���?             F@                                   �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  Pl@����>�?            �B@       	                           �?      �?             2@       
                        `ff�?�z�G��?             $@                                 �`@և���X�?             @                                   �?      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                      	             �?      �?              @        ������������������������       �                     �?                                ����?؇���X�?             @                                  `Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   `P@�}�+r��?
             3@       ������������������������       �        	             2@        ������������������������       �                     �?               2                    �?0� }��?�            �q@               %                   @m@r�q��?             B@               $                 ����?X�<ݚ�?             "@               #                    �?�q�q�?             @       !       "                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        &       -                   pc@�>����?             ;@       '       ,                    �? �q�q�?             8@        (       +                    �?�����H�?             "@       )       *                    �J@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        .       /                    �?�q�q�?             @        ������������������������       �                     �?        0       1                    _@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       ^                    �R@@�?��K�?�            �n@       4       7                    Z@��D�܇�?�            �n@        5       6                    @�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        8       ]                   �a@�1e�3��?�            �m@       9       :                    @J@p=
ףp�?d             d@        ������������������������       �        %            �O@        ;       N                    �?�Ι����??            @X@       <       G                   Pl@�Z��L��?.            �Q@       =       >                   Ph@����?�?            �F@       ������������������������       �                     @@        ?       @                    �?$�q-�?	             *@        ������������������������       �                     @        A       B                    �?�����H�?             "@        ������������������������       �                     @        C       D                 ����?r�q��?             @        ������������������������       �                     @        E       F                    @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        H       I                    Z@R�}e�.�?             :@        ������������������������       �                     "@        J       M                   (q@j���� �?             1@        K       L                 `ff�?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        O       \                    �?�θ�?             :@       P       [                   �`@�q�q�?             2@       Q       X                    �?      �?             (@       R       W                   �p@      �?             $@       S       V                   �Z@r�q��?             @        T       U                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        Y       Z                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        0             S@        _       `                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        b       g                    �?=&C��?6            �T@        c       d                   0n@��+7��?             7@       ������������������������       �                     ,@        e       f                    �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        h       u                   �b@z�G�z�?(             N@       i       p                    �?t��ճC�?              F@       j       k                   �`@ �q�q�?             8@       ������������������������       �                     1@        l       m                 ����?؇���X�?             @        ������������������������       �                     @        n       o                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        q       r                   `]@ףp=
�?             4@        ������������������������       �                     $@        s       t                    n@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        v       }                    �?     ��?             0@       w       x                   �\@�q�q�?             (@        ������������������������       �                     @        y       z                    @����X�?             @        ������������������������       �                     @        {       |                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               �                    �K@��&0n�?�            @t@       �       �                 033@(��6�ռ?�             k@       �       �                    �?�f�¦ζ?�            �j@       �       �                   Pd@@]����?n            @f@       �       �                    �I@0���ަ?k            �e@       �       �                    P@��d��?J             ^@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   `_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        G            @]@        �       �                    �?�1�`jg�?!            �K@       �       �                    �J@�&=�w��?            �J@        �       �                   �V@���}<S�?             7@        ������������������������       �                     �?        �       �                 ����?���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                     >@        �       �                   0f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0q@4?,R��?             B@       ������������������������       �                     9@        �       �                    �?�eP*L��?             &@       �       �                   pg@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��ɜ|��?B            �Z@       �       �                    �Q@�חF�P�?'             O@       �       �                    ]@���5��?$            �L@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@�NW���?"            �J@        �       �                    �?     ��?             0@       �       �                   �_@�r����?             .@        �       �                 @33�?���Q��?             @        ������������������������       �                      @        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        �       �       
             �?�?�|�?            �B@       ������������������������       �                     8@        �       �                   �c@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �Z@k��9�?            �F@        ������������������������       �                     @        �       �                    @O@D^��#��?            �D@       �       �                    �?�'�=z��?            �@@       �       �                    �?��}*_��?             ;@       �       �                   �i@������?	             1@       �       �                    @N@����X�?             ,@       �       �                   @g@r�q��?             (@       �       �                   �e@�<ݚ�?             "@       �       �                   �V@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���Q��?             $@        ������������������������       �                      @        �       �                    �L@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `ff @      �?              @       �       �                     P@؇���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  K�ۚ��?�)|�� �?�թX���?��թX��?
��֢P�?_�/���?F]t�E�?]t�E]�?۶m۶m�?�$I�$I�?      �?                      �?���L�?�u�)�Y�?      �?      �?333333�?ffffff�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?      �?                      �?              �?              �?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        (�����?�5��P�?              �?      �?        Տ3�ҵ�?�Y�EI�?UUUUUU�?�������?�q�q�?r�q��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?h/�����?�Kh/��?UUUUUU�?�������?�q�q�?�q�q�?UUUUUU�?�������?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ~*! 秲?�����?���Zeñ?�T���?UUUUUU�?UUUUUU�?              �?      �?        W'u_�?�/���?ffffff�?333333�?              �?���fy�?�Y�D�a�?��Vؼ?���.�d�?l�l��?��I��I�?              �?;�;��?�؉�؉�?              �?�q�q�?�q�q�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�;�;�?'vb'vb�?              �?ZZZZZZ�?�������?9��8���?�q�q�?      �?                      �?              �?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?      �?      �?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?              �?      �?        �����\�?�%���?zӛ����?Y�B��?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?t�E]t�?�E]t��?UUUUUU�?�������?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?�������?�������?              �?      �?              �?      �?�������?�������?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        <ݚ)�?����[�?�Tx*<�?��zX=��?��4>2��?�Ե��?�g<��?�as�Ü?�Z��D�?��4��g�?�������?�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        A��)A�?�־a�?tHM0���?�x+�R�?ӛ���7�?d!Y�B�?              �?�.�袋�?F]t�E�?      �?                      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �8��8��?r�q��?      �?        t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��G&�;�?�rp�_��?�Zk����?��RJ)��?�}��?��Gp�?      �?      �?      �?                      �?萚`���?�x+�R�?      �?      �?�������?�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?*�Y7�"�?к����?      �?        �؉�؉�?;�;��?      �?                      �?�������?333333�?              �?      �?        [�[��?�'}�'}�?              �?�]�ڕ��?,Q��+�?|��|�?|���?_B{	�%�?B{	�%��?xxxxxx�?�?�m۶m��?�$I�$I�?�������?UUUUUU�?9��8���?�q�q�?      �?      �?              �?      �?                      �?      �?                      �?      �?        �������?333333�?              �?      �?      �?      �?                      �?              �?      �?      �?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJc`>yhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         t                    �?.��X~��?�           ��@              9                    �?r٣����?�            �v@                                  @L@,Z0R�?�             m@                                  �?�d���?m            �e@                                  @G@�h����?i             e@        ������������������������       �        4            @T@                                ����?XB���?5            �U@                                  �?���7�?'            �P@        	       
                   �p@�C��2(�?             6@       ������������������������       �                     *@                                   f@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @                                   �?`���i��?             F@        ������������������������       �                     *@                      	             �?�g�y��?             ?@                                  �c@�����H�?             "@                                  �G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                     5@                                  `]@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @               4                 ����?>���Rp�?*             M@              3                    �?>a�����?$            �I@              *                   Hp@�:pΈ��?#             I@              )                    �?�L���?            �B@              $                    d@ףp=
�?             >@               !                    �Q@�nkK�?             7@       ������������������������       �                     5@        "       #                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       &                    �?����X�?             @       ������������������������       �                     @        '       (                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        +       .                    �M@�	j*D�?
             *@        ,       -                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        /       0                    `@      �?              @        ������������������������       �                     @        1       2                 ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        5       8                    �?؇���X�?             @       6       7                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        :       G                    �?���nU��?Y            ``@        ;       >                    �?��S�ۿ?             >@        <       =                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       F                    �? ��WV�?             :@       @       E                    V@���N8�?             5@        A       D                    @K@z�G�z�?             @        B       C                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     @        H       k                    �?&�����?D            @Y@       I       `                    �?     ��?6             T@       J       M                   �X@d��0u��?(             N@        K       L                    �J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        N       W                   Pb@�2����?%            �K@       O       R                   @E@�C��2(�?            �@@        P       Q                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        S       T                   p@XB���?             =@       ������������������������       �                     1@        U       V                   @^@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        X       _                   0m@���!pc�?             6@       Y       Z                   �e@և���X�?             ,@        ������������������������       �                     @        [       ^                    �F@�eP*L��?             &@        \       ]                   @b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        a       b                   �k@���Q��?             4@        ������������������������       �                     @        c       f                    �?�n_Y�K�?
             *@        d       e                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        g       h                    @F@      �?              @        ������������������������       �                     @        i       j                   �q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        l       o                   �Y@��s����?             5@        m       n                    �J@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        p       q                   �l@�IєX�?             1@       ������������������������       �        
             .@        r       s                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       �       	             �?�����?�            0w@       v       �                   �a@ ~�����?�            �u@       w       �                    �P@��u���?�            pp@       x       }                    �?��*;�?�             n@        y       z                   (s@@4և���?             E@       ������������������������       �                     C@        {       |                   @[@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                    �? ���v��?}            �h@               �                    �H@�z�G��?             4@        ������������������������       �                     @        �       �                 ����?���Q��?
             .@        ������������������������       �                      @        �       �                    �?��
ц��?             *@       �       �                    a@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�x�E~�?p            @f@        ������������������������       �                     E@        �       �                 033@г�wY;�?U             a@       �       �                    �?P����?J            �]@        ������������������������       �                     C@        �       �                 hff�?�(\����?-             T@        �       �                    _@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @i@`׀�:M�?*            �R@        �       �                   `_@(;L]n�?             >@       ������������������������       �                     ;@        �       �                    Y@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     F@        �       �                   �\@�����H�?             2@        �       �                    �J@z�G�z�?             $@        �       �                    @J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�㙢�c�?             7@       �       �                    _@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                   �[@���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �N@���R�?4            @T@       �       �                    @&����?*            @P@       �       �                    h@Ȩ�I��?#            �J@        ������������������������       �        	             .@        �       �                    �?p�ݯ��?             C@       �       �                    @M@j���� �?             A@       �       �       
             �?      �?             :@        �       �                    �?8�Z$���?	             *@        �       �                   Pb@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �r@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    @H@8�Z$���?	             *@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                   @l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0n@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �       
             �?      �?
             0@       �       �                    �?�����H�?             "@       �       �                   pc@r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             ;@       �       �                    �L@؇���X�?             5@       �       �                    c@�IєX�?             1@        �       �                   �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 `ff�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  ��� ���?���o���?>���>�?|���?�FX�i��?	�=��ܳ?�:���C�?Ȥx�L��?۶m۶m�?�$I�$I�?      �?        GX�i���?�{a���?�.�袋�?F]t�E�?]t�E�?F]t�E�?      �?        9��8���?�q�q�?      �?                      �?F]t�E�?F]t�E�?      �?        ��{���?�B!��?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?              �?        �������?UUUUUU�?              �?      �?        �i��F�?GX�i���?�������?�?��Q���?�Q����?}���g�?L�Ϻ��?�������?�������?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?                      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        vb'vb'�?;�;��?�������?333333�?      �?                      �?      �?      �?      �?        �������?�������?              �?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?T���0��?V���g�?�?�������?      �?      �?              �?      �?        ;�;��?O��N���?�a�a�?��y��y�?�������?�������?      �?      �?      �?                      �?              �?              �?              �?� w�l��?�&��?      �?      �?�?�������?�������?�������?      �?                      �?��7�}��?� O	��?]t�E�?F]t�E�?      �?      �?      �?                      �?GX�i���?�{a���?      �?        UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?        ]t�E�?t�E]t�?�������?UUUUUU�?      �?                      �?              �?      �?        �������?333333�?              �?;�;��?ى�؉��?�������?�������?      �?                      �?      �?      �?              �?�������?�������?      �?                      �?�a�a�?z��y���?      �?      �?      �?                      �?�?�?              �?      �?      �?      �?                      �?|?��o��?!��d�?A_���?�}A_�?��2�*��?J�y�z��?�������?DDDDDD�?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        1ogH�۩?�y;Cb�?333333�?ffffff�?              �?�������?333333�?              �?�؉�؉�?�;�;�?333333�?�������?      �?                      �?              �?p�\��?����G�?              �?�?�?'u_[�?�V'u�?              �?�������?333333�?UUUUUU�?�������?              �?      �?        к����?��L��?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?�q�q�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?d!Y�B�?�7��Mo�?�q�q�?��8��8�?      �?                      �?333333�?�������?              �?      �?      �?      �?                      �?��ӭ�a�?�)O�?�����?�����?�	�[���?+�R��?              �?Cy�5��?^Cy�5�?ZZZZZZ�?�������?      �?      �?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        ;�;��?;�;��?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?              �?      �?      �?�q�q�?�q�q�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?�?�?�������?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJا�LhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKͅ�h��B@3         �       	             �?znt��s�?�           ��@              q                    �?�4�س�?v           ��@              \       
             �?��ɉ�?�            `x@                                  �?<
ףp-�?�             t@               
                    �?��Q��?             4@              	                    �?"pc�
�?             &@                                   �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   `@X�<ݚ�?             "@                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   p@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               %                    �?ףp=
�?�            �r@               "                   �e@�+Ĺ+�?3            �T@                               ����?P���Q�?1             T@        ������������������������       �                    �A@                                   �?�:�^���?            �F@                                  �?�7��?            �C@                                 pc@ ��WV�?             :@       ������������������������       �                     8@                                   �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �h@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?                !                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        #       $                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        &       [                    �R@T���.�?�             k@       '       J                 ����?��f��?�            �j@       (       3                    �?؇���X�?K            �]@        )       .                   `a@8����?             7@        *       +                   �n@�q�q�?             "@        ������������������������       �                     @        ,       -                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        /       2                   pl@@4և���?             ,@        0       1                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        4       I                     P@8��8���?>             X@       5       <                    @K@�?�'�@�?3             S@       6       ;                    �?P���Q�?             D@       7       8                    �?�>����?             ;@       ������������������������       �                     8@        9       :                    r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@        =       >                   0h@�<ݚ�?             B@       ������������������������       �                     3@        ?       F                    @M@��.k���?
             1@       @       A                    W@���Q��?             $@        ������������������������       �                      @        B       C                   �`@      �?              @        ������������������������       �                     @        D       E                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        G       H                 433�?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     4@        K       P                     G@��s��?9            �W@        L       O                    �?"pc�
�?             &@       M       N                     F@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        Q       Z                    �?�Ń��̧?3             U@       R       W                   �_@(;L]n�?&             N@        S       T                   �^@ףp=
�?             $@       ������������������������       �                      @        U       V                   po@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        X       Y                    c@p���?              I@       ������������������������       �                    �H@        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     @        ]       p                   �r@���L��?,            �Q@       ^       e                   ph@�����D�?*            @P@        _       `                    �F@�FVQ&�?            �@@        ������������������������       �                     �?        a       b                    a@      �?             @@       ������������������������       �                     ;@        c       d                   @e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        f       o                   �n@     ��?             @@       g       h                    �?\X��t�?             7@        ������������������������       �                     @        i       j                     F@�E��ӭ�?             2@        ������������������������       �                     @        k       n                    @N@�r����?
             .@       l       m                   pm@@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        r       �                 ����?��"�ű�?�            �i@       s       �                    �?T&ss��?]            �`@       t       }                   `]@L�'�7��?P            @]@        u       v                    �?>���Rp�?             =@        ������������������������       �                     &@        w       |                    �?b�2�tk�?             2@       x       y                   @b@������?             .@        ������������������������       �                      @        z       {                   @f@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ~       �                   Pb@���7�?=             V@              �                    �?�g<a�?6            @S@        ������������������������       �                    �A@        �       �                   �r@���N8�?             E@       �       �                 ����? ���J��?            �C@       ������������������������       �                     @@        �       �                 833�?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@       �       �                    j@ףp=
�?             $@        �       �                    �N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?X�<ݚ�?             2@        ������������������������       �                     @        �       �                    �?և���X�?
             ,@        ������������������������       �                     �?        �       �                     M@�n_Y�K�?	             *@       �       �                   @`@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�xGZ���?&            �Q@       �       �                   @l@��]�T��?            �D@        �       �                    �?z�G�z�?	             .@       �       �                    �?d}h���?             ,@        ������������������������       �                      @        �       �                     L@      �?             @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 033@ȵHPS!�?             :@       �       �                    �M@HP�s��?             9@        ������������������������       �                     $@        �       �                    �?�r����?             .@        ������������������������       �                     $@        �       �                   `a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �_@V�a�� �?             =@        ������������������������       �                     1@        �       �                   �`@      �?
             (@        �       �                   �r@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����X�?             @        ������������������������       �                      @        �       �                   �e@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?~=�r�?[            `a@        �       �                   �o@���>4��?             <@       �       �                   �`@     ��?             0@       �       �                    �L@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �                   @g@�g+��@�?G            �[@       �       �                    �? '��h�?F            @[@        ������������������������       �                     F@        �       �                    @L@$�q-�?+            @P@       ������������������������       �        %             J@        �       �                 ����?�n_Y�K�?             *@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ����?��}t��?�L��L��?��"��"�?�����?�����?�������?�����L�?ffffff�?�������?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?r�q��?�q�q�?      �?      �?      �?                      �?�������?333333�?      �?                      �?�������?�������?���ˊ��?(፦ί�?�������?ffffff�?              �?l�l��?}�'}�'�?�A�A�?��[��[�?;�;��?O��N���?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�@q�8P�?�����u�?��XQ�?A�Ե��?�$I�$I�?۶m۶m�?8��Moz�?d!Y�B�?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?      �?        �$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?�������?�������?y�5���?������?�������?ffffff�?h/�����?�Kh/��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?9��8���?              �?�?�������?333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?      �?                      �?              �?�X�0Ҏ�?q�����?F]t�E�?/�袋.�?�������?�������?              �?      �?                      �?�a�a�?��<��<�?�?�������?�������?�������?              �?      �?      �?              �?      �?        {�G�z�?\���(\�?              �?      �?                      �?      �?        _�_��?��:��:�?z�z��?z�z��?|���?>����?      �?              �?      �?              �?�������?�������?              �?      �?              �?      �?��Moz��?!Y�B�?      �?        r�q��?�q�q�?      �?        �?�������?�$I�$I�?n۶m۶�?              �?      �?              �?                      �?      �?        ��q9�?�Ѹ���?�)F�?= Y���?�������?���?�i��F�?GX�i���?      �?        �8��8��?9��8���?wwwwww�?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?                      �?�.�袋�?F]t�E�?���8+�?�cj`?      �?        ��y��y�?�a�a�?��-��-�?�A�A�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?/�袋.�?F]t�E�?�������?�������?�������?�������?              �?      �?              �?                      �?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?        ى�؉��?;�;��?�m۶m��?�$I�$I�?              �?      �?                      �?�A�A�?�_�_�?KԮD�J�?jW�v%j�?�������?�������?۶m۶m�?I�$I�$�?              �?      �?      �?      �?      �?              �?      �?                      �?              �?��N��N�?�؉�؉�?q=
ףp�?{�G�z�?      �?        �������?�?      �?        333333�?�������?      �?                      �?              �?a���{�?��{a�?              �?      �?      �?�������?�������?      �?                      �?�$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?        gXp�l��?c�>ZMB�?n۶m۶�?I�$I�$�?      �?      �?]t�E�?F]t�E�?      �?                      �?�������?�������?      �?                      �?UUUUUU�?�������?      �?                      �?���+c��?Nq��$�?���]8��?�w� z|�?      �?        �؉�؉�?;�;��?      �?        ;�;��?ى�؉��?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�|MhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK녔h��B�:         �                    �?�ܲ�}��?�           ��@              Q                    �? �*�bf�?           �z@              ,                    �?^ex�Ñ�?�             q@              )                 ���@p���p�?�            �i@              &                   �g@8?W���?}             i@                                 pl@�Q �?{            �h@                                  �?`�LVXz�?>            �X@       ������������������������       �        9            �W@        	                           �?z�G�z�?             @       
                           @L@      �?             @        ������������������������       �                      @                                  `b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   �?������?=            @X@        ������������������������       �                      @                                   �?�KM�]�?<            �W@        ������������������������       �                     9@               %                    �?؇���X�?(            �Q@                                  @L@6YE�t�?%            �P@                                 �n@�&=�w��?            �J@                      	             �?r�q��?             (@                                  �\@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �D@                                    �?�n_Y�K�?             *@                                @33�?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        !       "       	             �?X�<ݚ�?             "@        ������������������������       �                     �?        #       $                   �_@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        '       (                    �D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        *       +                   �]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        -       B                   `_@�v:���?/             Q@       .       A                    �?��Zy�?            �C@       /       @                    _@��
P��?            �A@       0       ;                 ����?��>4և�?             <@       1       :                   `]@�d�����?             3@       2       3                   @[@�eP*L��?	             &@        ������������������������       �                     @        4       9                 ����?      �?              @       5       8                    �?����X�?             @       6       7                    @F@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        <       ?                    �?�q�q�?             "@        =       >                    `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        C       N                    �?ܷ��?��?             =@       D       I                   �i@�>����?             ;@        E       H                 @33�?r�q��?             @       F       G                   h@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        J       K                   d@���N8�?             5@       ������������������������       �        
             .@        L       M                   @c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        O       P                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       S                   �\@x�(�3��?a            @c@        ������������������������       �                    �A@        T       �                    �?�n\�GZ�?J            �]@       U       �                    �Q@\X��t�?:             W@       V       q                    �?�&!��?8            �U@       W       p                   �d@�F�j��?             �J@       X       i                 `ff�?�zv�X�?             F@       Y       d                    �?X�<ݚ�?             ;@       Z       c                 `ff�?�q�q�?             (@       [       \                   �\@���!pc�?
             &@        ������������������������       �                     @        ]       b                   0a@և���X�?             @       ^       a                   �_@      �?             @        _       `                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        e       f                    �?������?             .@        ������������������������       �                     "@        g       h                    �G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        j       o                   0b@�t����?             1@        k       l       
             �?���Q��?             @        ������������������������       �                     �?        m       n                   pj@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     "@        r       {                    �?r٣����?            �@@        s       t                    @L@X�<ݚ�?             "@        ������������������������       �                      @        u       z                    �?����X�?             @       v       w                   xu@r�q��?             @       ������������������������       �                     @        x       y                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        |       �                   �e@r�q��?             8@       }       �                    n@�C��2(�?             6@       ~                           @K@؇���X�?
             ,@       ������������������������       �                      @        �       �                    �N@�q�q�?             @       �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�<ݚ�?             ;@        �       �                    @O@��
ц��?             *@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                 ����?��z�}T�?�             s@        �       �                    �?���Q��?.            �R@        �       �                    �?����>�?            �B@        ������������������������       �                     *@        �       �                    �?�q�q�?             8@       �       �                    h@�E��ӭ�?	             2@        ������������������������       �                     @        �       �                   @`@�r����?             .@        �       �                    _@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                   �]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�˹�m��?             C@       ������������������������       �                     ;@        �       �                 @33�?���!pc�?             &@       �       �                     I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��0���?�            �l@       �       �                   P`@x�}b~|�?�            �l@       �       �                    �?��w#'�?e            `d@       �       �                    �?Ц�f*�?E            �[@        �       �                    @H@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?p� V�?A            �Y@       �       �                   `_@�Fǌ��?/            �S@       ������������������������       �        &            �M@        �       �                   �j@P���Q�?	             4@        �       �                    �J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   `c@ �q�q�?             8@       ������������������������       �                     3@        �       �                    �?z�G�z�?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? �h�7W�?             �J@        �       �                     N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0p@p���?             I@       ������������������������       �                    �B@        �       �                   �_@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                     O@&����?+            @P@       �       �                   �V@^(��I�?&            �K@        ������������������������       �                      @        �       �                    �?�T`�[k�?%            �J@        �       �                     E@���Q��?             @        ������������������������       �                     �?        �       �                   `c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �M@     ��?              H@       �       �                    �?      �?             D@       �       �                    l@$�q-�?             :@        ������������������������       �                     (@        �       �                    �?؇���X�?             ,@        ������������������������       �                     @        �       �                   �n@z�G�z�?	             $@        ������������������������       �                     �?        �       �                    q@�����H�?             "@        ������������������������       �                     @        �       �                    c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?d}h���?             ,@       �       �                     H@      �?             (@        ������������������������       �                      @        �       �                     M@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    b@      �?              @       �       �                   �Y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �t�b��#     h�h)h,K ��h.��R�(KK�KK��hi�B�  ����u��?/�E��?�B�(���?z�����?ZP�9���?��J��?�E|���?C��ڸ?F��s�?�����`�?x9/���??4և���?�~�@��?[�R�֯�?      �?        �������?�������?      �?      �?      �?              �?      �?              �?      �?              �?        |q���
�? tT����?              �?�k(���?(�����?      �?        ۶m۶m�?�$I�$I�?'�l��&�?e�M6�d�?tHM0���?�x+�R�?�������?UUUUUU�?333333�?�������?              �?      �?              �?              �?        ى�؉��?;�;��?      �?      �?              �?      �?        �q�q�?r�q��?      �?              �?      �?              �?      �?              �?        �������?333333�?      �?                      �?�������?�������?      �?                      �?<<<<<<�?�������?\��[���?� � �?_�_��?PuPu�?۶m۶m�?I�$I�$�?Cy�5��?y�5���?t�E]t�?]t�E�?      �?              �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?              �?��=���?a���{�?�Kh/��?h/�����?�������?UUUUUU�?�������?�������?      �?                      �?      �?        ��y��y�?�a�a�?      �?        �������?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�wL��?(�Y�	q�?              �?�O��O��?4X�3X��?��Moz��?!Y�B�?S֔5eM�?֔5eMY�?:�&oe�?��sHM�?�袋.��?��.���?r�q��?�q�q�?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?        wwwwww�?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�?<<<<<<�?�������?333333�?              �?      �?      �?              �?      �?                      �?      �?        |���?>���>�?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        UUUUUU�?�������?F]t�E�?]t�E�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?              �?        �q�q�?9��8���?�؉�؉�?�;�;�?              �?      �?                      �?ր+ր+�?�u�u�?�������?333333�?�u�)�Y�?���L�?      �?        �������?�������?�q�q�?r�q��?              �?�������?�?      �?      �?      �?                      �?      �?        UUUUUU�?�������?              �?�������?�������?      �?                      �?^Cy�5�?��P^Cy�?              �?t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?      �?        ��e�:}�?cAs�X��?Lg1��t�?�YLg1�?��\w�آ?f5�8t��?�־a�?!O	� �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?��,�?����`�?�3���?1���M��?              �?�������?ffffff�?�������?�������?              �?      �?                      �?UUUUUU�?�������?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?"5�x+��?��sHM0�?UUUUUU�?UUUUUU�?              �?      �?        {�G�z�?\���(\�?              �?;�;��?�؉�؉�?      �?                      �?�����?�����?J��yJ�?�7�}���?      �?        "5�x+��?���!5��?333333�?�������?              �?      �?      �?      �?                      �?      �?      �?      �?      �?;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?        �q�q�?�q�q�?              �?�������?�������?              �?      �?        ۶m۶m�?I�$I�$�?      �?      �?      �?        �������?�������?              �?      �?                      �?      �?      �?�������?�������?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�#vhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         �                    �?���-�g�?�           ��@                                  f@(�f����?	           �z@                                   �?����?Q            @`@                                 @e@����1�?-            @R@                                 �]@p��%���?+            @Q@        ������������������������       �                     ?@                                   �?�KM�]�?             C@               	                    �D@      �?             @        ������������������������       �                     �?        
                           �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   �?�IєX�?             A@                                   �?���Q��?             @        ������������������������       �                     �?                                  �U@      �?             @                                 `Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        $            �L@               W                   �a@��Xd���?�            �r@              V                    �R@(L���?            �j@              A                   ``@��?��:�?~            �j@               @                    �?���Fi�?6            �T@              +                    `@�iޤ��?-            �P@                                   �?� ��1�?            �D@        ������������������������       �                     @        !       *                    �L@������?            �B@       "       )                    @L@z�G�z�?             4@       #       $                    g@�����H�?             2@        ������������������������       �                     �?        %       &                   (p@�IєX�?             1@       ������������������������       �        
             $@        '       (                   `p@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        ,       3                    �?��
ц��?             :@        -       2                    �?�����H�?             "@       .       /                   �l@      �?              @        ������������������������       �                     @        0       1                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        4       5                    �K@������?             1@        ������������������������       �                      @        6       ?                    t@X�<ݚ�?             "@       7       >                   �s@և���X�?             @       8       =                   `n@���Q��?             @       9       <                    �?�q�q�?             @       :       ;                   @k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@        B       U                   pn@����?H            @`@        C       P                   0`@(2��R�?             �M@       D       O       
             �?      �?             H@       E       H                    �K@�#-���?            �A@        F       G                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        I       N                    �?h�����?             <@        J       K                    �?؇���X�?             @       ������������������������       �                     @        L       M                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             5@        ������������������������       �                     *@        Q       T                   pb@�eP*L��?             &@       R       S       	             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        (            �Q@        ������������������������       �                      @        X       �                   0f@yÏP�?9            �T@       Y       r                   �o@���L��?5            �S@       Z       o       	             �?�q�q�?             E@       [       n                   n@     ��?             @@       \       a                    �?J�8���?             =@        ]       `                    �?8�Z$���?             *@       ^       _                    @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        b       c                   �g@      �?             0@        ������������������������       �                     @        d       e                     D@�n_Y�K�?	             *@        ������������������������       �                     �?        f       g                 hff�?�q�q�?             (@        ������������������������       �                     @        h       i                   @b@�q�q�?             @        ������������������������       �                     �?        j       m                   �l@z�G�z�?             @        k       l                     K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        p       q                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        s       �                    �?�8��8��?             B@        t       u                    �?z�G�z�?             .@        ������������������������       �                     �?        v                           �?؇���X�?
             ,@       w       ~                    �?z�G�z�?             $@       x       }                   �z@�<ݚ�?             "@       y       |                 `ff�?      �?              @        z       {                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                     @        �       �                    �?���
.��?�            0s@       �       �                   h@(���h�?�            �i@       �       �                   �c@`n31�=�?�            `i@       �       �       	             �?�nkK�?w             g@        �       �                 ���@dP-���?9            �W@       �       �                   �t@0�>���?7            �V@       �       �       
             �?`Ӹ����?6            �V@        �       �                   h@"pc�
�?             &@       ������������������������       �                     @        �       �                   @]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �G@pY���D�?1            �S@        �       �                    �?@4և���?             <@        ������������������������       �                      @        �       �                   0n@ףp=
�?             4@       ������������������������       �        	             *@        �       �                    �F@����X�?             @        ������������������������       �                     @        �       �                   �]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �I@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        >            �V@        �       �                     R@�S����?
             3@       ������������������������       �        	             0@        ������������������������       �                     @        ������������������������       �                      @        �       �                 ����?4�M�f��??            �Y@       �       �                    �?��paR�?,             Q@       �       �                    �?�q�q�?              H@       �       �                    @D@8�Z$���?            �C@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�#-���?            �A@       �       �                    �?�g�y��?             ?@        �       �                   @_@      �?             0@       �       �                   @[@      �?              @        �       �                 @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        �       �                   �c@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �c@X�<ݚ�?             "@       �       �                   �a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �p@�G�z��?             4@        �       �                    �?�z�G��?             $@        ������������������������       �                      @        �       �                   �f@      �?              @       �       �                    @I@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �r@z�G�z�?             $@        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    @M@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 033�?@�0�!��?             A@       �       �                    a@ףp=
�?             >@       �       �                    �?     ��?	             0@        �       �                   0p@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     ,@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  lk�w��?J��	.�?�a�H��?�':ݭ��?�����?n�Fn�F�?Ĉ#F��?�Ν;w��?ہ�v`��?�g��%�?              �?(�����?�k(���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�?�������?333333�?      �?              �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?                      �? cţr�?8�W#��?w�qG��?⎸#��?��χ��?����?��FS���?�C.+J�?�rv��?��Dz�r�?������?������?      �?        к����?��g�`��?�������?�������?�q�q�?�q�q�?      �?        �?�?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?�؉�؉�?�;�;�?�q�q�?�q�q�?      �?      �?      �?              �?      �?      �?                      �?      �?        �?xxxxxx�?              �?�q�q�?r�q��?�$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?                      �?              �? �����?~�~��?'u_[�?=�"h8��?      �?      �?_�_�?�A�A�?�$I�$I�?�m۶m��?      �?                      �?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?              �?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?      �?              �?                      �?      �?        Q��+Q�?W�v%jW�?��o��o�?�4H�4H�?UUUUUU�?UUUUUU�?      �?      �?�rO#,��?|a���?;�;��?;�;��?333333�?�������?      �?                      �?      �?              �?      �?              �?;�;��?ى�؉��?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?              �?              �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?        �$I�$I�?۶m۶m�?�������?�������?�q�q�?9��8���?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?              �?              �?      �?        �}�?��F���?��߁��?<��;�?J��8D�?Ztl��?�Mozӛ�?d!Y�B�?�����F�?W�+�ɵ?��=��=�?�!�!�??�>��?l�l��?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?a~W��0�?�3���?n۶m۶�?�$I�$I�?      �?        �������?�������?      �?        �m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?              �?      �?        (������?^Cy�5�?      �?                      �?              �?�������?�������?�?�������?UUUUUU�?�������?;�;��?;�;��?      �?      �?      �?                      �?�A�A�?_�_�?��{���?�B!��?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?              �?              �?      �?      �?                      �?r�q��?�q�q�?�������?UUUUUU�?              �?      �?                      �?�������?�������?ffffff�?333333�?      �?              �?      �?�������?333333�?              �?      �?              �?        �������?�������?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?�������?ZZZZZZ�?�������?�������?      �?      �?۶m۶m�?�$I�$I�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ>hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�7         v                    �?
���P��?�           ��@              O                    �?��I�C�?�            @x@              2                    �?��y*�?�            r@              /                 ���@�L�3�?�            �k@              .                   �g@��$xtW�?�            �j@              	                   �O@ �h�7W�?�            �j@                                   `Q@      �?              @       ������������������������       �                     @        ������������������������       �                     @        
       -                   e@ =[y��?}            �i@                                  @L@�IєX�?]             c@                                 �d@@�n�1�?I            @_@                                 �b@��d��?G             ^@       ������������������������       �        +            @Q@                      
             �?���J��?            �I@       ������������������������       �                     9@                                   @H@ ��WV�?             :@                                  c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@                                   �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?               ,                    �?      �?             <@              '       	             �?�q�q�?             8@                                   �?ҳ�wY;�?             1@                                  �O@z�G�z�?             $@        ������������������������       �                     @                                   �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        !       &                    �?և���X�?             @       "       %                    �?���Q��?             @       #       $                    @N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        (       )                   �?؇���X�?             @       ������������������������       �                     @        *       +                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �I@        ������������������������       �                     �?        0       1       
             �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        3       L                    �?4�	~���?.            @Q@       4       E                    �?��mo*�?%            �M@       5       6                    �?�����H�?            �F@        ������������������������       �                     (@        7       D                    �?6YE�t�?            �@@       8       C                    @N@r�q��?             >@       9       @                   �d@\-��p�?             =@       :       ;                 @33�?$�q-�?             :@       ������������������������       �                     5@        <       ?                 @33�?���Q��?             @       =       >                    `@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        A       B                   `m@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        F       G                   �_@X�Cc�?	             ,@        ������������������������       �                     @        H       K                    �?      �?              @       I       J                    s@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        M       N                   `@z�G�z�?	             $@       ������������������������       �                      @        ������������������������       �                      @        P       m                   �b@�I{A�?;            �X@       Q       X                 ����?�=A�F�?.             S@        R       U                    �?���Q��?             $@       S       T                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        V       W                    �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        Y       l       	             �?��2(&�?(            �P@       Z       a                    �?�?�<��?'            @P@       [       \                   �r@P�Lt�<�?             C@       ������������������������       �                     A@        ]       `                   �_@      �?             @       ^       _                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        b       c                    �?������?             ;@        ������������������������       �                      @        d       i                    c@z�G�z�?             9@       e       f                 033�?؇���X�?
             5@       ������������������������       �                     1@        g       h                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        j       k                    @M@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        n       u                    `@�LQ�1	�?             7@        o       t                    �?      �?              @       p       q                    �?����X�?             @        ������������������������       �                     @        r       s       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        w       �                   �b@H~4o]�?�            �u@       x                          @f@�C��2(�?�            0q@        y       ~                    �?@��,B�?8            �V@        z       }                    �?P���Q�?             4@        {       |                   �\@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     "@        ������������������������       �        ,            �Q@        �       �                    �?�LQ�1	�?p             g@        �       �                   �_@R�}e�.�?             :@        �       �                    @N@�q�q�?             (@       �       �                   �r@      �?              @       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �       	             �?؇���X�?
             ,@       �       �                   �`@$�q-�?	             *@        �       �                    �J@r�q��?             @        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   p`@���1���?`            �c@       �       �                    �?���l��?C            �[@       �       �                    @L@�(�Tw�?/            �S@       ������������������������       �                     D@        �       �                   @i@P�Lt�<�?             C@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?�'�`d�?            �@@        �       �                    �?��Q��?
             4@        ������������������������       �                     @        �       �                    @��S���?             .@       �       �                   q@��
ц��?             *@       �       �                    `@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             *@        �       �                    �?��k=.��?            �G@        �       �                    @E@ҳ�wY;�?
             1@        ������������������������       �                      @        �       �                    �?������?	             .@       ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        �       �                     P@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             >@       �       �                    @L@�nkK�?             7@       ������������������������       �        	             0@        �       �                   pb@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����X�?             @        �       �                   �j@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?R_u^|�?*            �Q@       �       �                    �?��<b���?             G@       �       �                    �?8^s]e�?             =@       �       �                   �p@��X��?             <@       �       �                 033�?      �?             8@       �       �                    @C@��
ц��?	             *@        ������������������������       �                     @        �       �                    �?���Q��?             $@        �       �                   d@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �                   0d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                     E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    _@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �                     0@        �       �                   �g@�J�4�?             9@        ������������������������       �                      @        �       �                    @���}<S�?             7@       �       �                   �p@���7�?             6@       ������������������������       �        	             2@        �       �                    �?      �?             @       �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  փmM���?>IY�8�??��W�?�/�~�Q�?:߄*�u�?��U�(�?=%�S�<�?־a��?����?��n�?�?��sHM0�?"5�x+��?      �?      �?      �?                      �?�������?�������?�?�?�rh��|�?����Mb�?�������?�?      �?        ______�?�?      �?        O��N���?;�;��?۶m۶m�?�$I�$I�?              �?      �?              �?        �������?�������?      �?                      �?      �?      �?�������?�������?�������?�������?�������?�������?      �?        333333�?�������?      �?                      �?۶m۶m�?�$I�$I�?333333�?�������?      �?      �?              �?      �?              �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?�$I�$I�?۶m۶m�?      �?                      �?];0���?F��Q�g�?�<�"h�?W'u_�?�q�q�?�q�q�?      �?        '�l��&�?e�M6�d�?�������?UUUUUU�?a����?�{a���?�؉�؉�?;�;��?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �m۶m��?%I�$I��?              �?      �?      �?�m۶m��?�$I�$I�?      �?                      �?              �?�������?�������?              �?      �?        K�Z�R��?[�R�֯�?6��P^C�?��k(��?333333�?�������?�������?UUUUUU�?      �?                      �?      �?      �?              �?      �?        t�E]t�?��.���? �����?�����?(�����?���k(�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?{	�%���?B{	�%��?      �?        �������?�������?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?              �?        ��Moz��?Y�B��?      �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        +���}��?5�� ��?F]t�E�?]t�E�?h�h��?`��_���?�������?ffffff�?F]t�E�?]t�E�?      �?                      �?              �?              �?Y�B��?��Moz��?�;�;�?'vb'vb�?�������?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?      �?        7a~W��?�3���?5'��Ps�?��蕱�?�A�A�?p��o���?              �?(�����?���k(�?      �?      �?              �?      �?                      �?'�l��&�?6�d�M6�?ffffff�?�������?              �?�������?�?�;�;�?�؉�؉�?ffffff�?333333�?      �?                      �?              �?              �?              �?br1���?g���Q��?�������?�������?      �?        �?wwwwww�?              �?�q�q�?r�q��?�������?�������?      �?                      �?              �?�������?�������?d!Y�B�?�Mozӛ�?              �?�$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?2~�ԓ��?�@�6�?��Moz��?��,d!�?	�=����?|a���?%I�$I��?n۶m۶�?      �?      �?�؉�؉�?�;�;�?              �?333333�?�������?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?      �?      �?      �?                      �?      �?                      �?      �?      �?              �?      �?                      �?�?�?      �?                      �?�z�G��?{�G�z�?              �?ӛ���7�?d!Y�B�?�.�袋�?F]t�E�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���GhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��B@6         R                    �?�/� d:�?�           ��@               +                 ����?V�lf��?�            �s@                                  �?�$
��
�?�            `j@                                   �?��Q��?             D@                                   Q@V������?            �B@                                 @a@��R[s�?            �A@                                  �?և���X�?             5@              	                    b@�q�q�?             (@        ������������������������       �                     @        
                          �p@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                  @^@�<ݚ�?             "@       ������������������������       �                     @                                  �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �                      @        ������������������������       �                     @                                  �O@�����?r            `e@                                   �P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  @n@ Df@��?n            �d@       ������������������������       �        :            �V@               *                   �g@�}�+r��?4             S@                                 �n@�?�|�?3            �R@                                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                !                   �?�k~X��?1             R@       ������������������������       �        +            @P@        "       )                    �?؇���X�?             @       #       $                    �?      �?             @        ������������������������       �                     �?        %       &                   @a@�q�q�?             @        ������������������������       �                     �?        '       (                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ,       3                    �?<W#.m��?E            @Z@        -       .                    �?��� ��?             ?@        ������������������������       �        	             ,@        /       2                    \@������?
             1@        0       1                    �L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        4       5                   �_@^��4m�?2            �R@        ������������������������       �                     9@        6       M                   Pe@`�(c�?!            �H@       7       @                   �j@�>$�*��?            �D@        8       9                 033�?�q�q�?             5@       ������������������������       �                     (@        :       ?                 ���@�<ݚ�?             "@       ;       >                    �?����X�?             @       <       =                   @a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        A       D                    �?z�G�z�?             4@        B       C                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        E       F                 `ff�?      �?             0@        ������������������������       �                     @        G       L       
             �?�����H�?             "@       H       I                    �?؇���X�?             @        ������������������������       �                     @        J       K                    �K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        N       Q                    �E@      �?              @        O       P                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        S       �                    @N@�X!���?            z@       T       �                    �?B`�I��?�            `r@        U       �                 ����?v�\!L^�?N            @^@       V       w                    �?�'�=z��?B            �X@       W       X                    �?>���Rp�?(             M@        ������������������������       �                     "@        Y       b                    T@����X�?!            �H@        Z       [                    �?���!pc�?             &@        ������������������������       �                     @        \       ]                    �և���X�?             @        ������������������������       �                     �?        ^       a                 @33�?      �?             @       _       `                    @D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        c       r                   �_@�S����?             C@        d       e                     E@�t����?             1@        ������������������������       �                     �?        f       m                    �?      �?
             0@        g       l                    �?؇���X�?             @       h       k                    �J@z�G�z�?             @       i       j                   `]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        n       q                   @f@�q�q�?             "@       o       p                   pn@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        s       t                   �b@���N8�?             5@       ������������������������       �                     3@        u       v                   po@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       y                   `g@��r._�?            �D@        ������������������������       �                     4@        z       {                   @h@�q�q�?             5@        ������������������������       �                     �?        |       }                    �?�z�G��?             4@       ������������������������       �                     $@        ~       �                    �M@���Q��?             $@              �                   �b@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���7�?             6@        �       �                    �F@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                    �?E�Vl��?m            �e@       �       �                    �?Xș���?S            �`@       �       �                    a@��(�?H            @\@       �       �                 ����?���1j	�?7            �U@       �       �                    �?ףp=
�?             I@       �       �                   �[@,���i�?            �D@        ������������������������       �                      @        �       �                    @L@$�q-�?            �C@       �       �                    �I@Pa�	�?            �@@        �       �                    �?��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �        
             2@        �       �                 ����?�q�q�?             @       �       �                   �Z@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     B@        �       �                    �?l��
I��?             ;@        ������������������������       �                     �?        �       �                   �a@R�}e�.�?             :@        �       �                   �a@X�<ݚ�?             "@       �       �                    �?և���X�?             @       �       �                    �K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   `q@�t����?             1@       �       �                   0c@�<ݚ�?             "@       �       �                 033@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�eP*L��?             6@       �       �                   ht@�G��l��?
             5@       �       �                 ����?D�n�3�?	             3@       �       �                   pf@     ��?             0@       �       �                    b@d}h���?             ,@       �       �                   �`@�8��8��?             (@        �       �                   @d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?P�Lt�<�?             C@        ������������������������       �                     �?        ������������������������       �                    �B@        �       �                    �?`Jj��?J             _@       �       �                    �?@3����?>             [@       �       �                   �a@      �?$             P@       �       �                    �?�X�<ݺ?             B@       �       �                 ����?�C��2(�?             6@        �       �                   �a@      �?              @       �       �                 `ff�?؇���X�?             @        ������������������������       �                     @        �       �                   `]@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �        	             ,@        ������������������������       �                     <@        ������������������������       �                     F@        �       �                    �?      �?             0@       �       �                     P@"pc�
�?             &@       �       �                   �V@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 hff�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  b�UK��?�U�)|�?�M�����?ud�@T:�?=:�oL�??�A��?ffffff�?�������?o0E>��?�g�`�|�?PuPu�?X|�W|��?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        ��w�?�A|�?�������?�������?      �?                      �?c��7�:�?��k���?      �?        �5��P�?(�����?*�Y7�"�?к����?      �?      �?      �?                      �?�8��8��?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?��	��	�?�����?�{����?�B!��?      �?        xxxxxx�?�?�������?�������?      �?                      �?      �?        �S�n�?�|����?              �?4և����?������?�����?�18���?UUUUUU�?UUUUUU�?      �?        �q�q�?9��8���?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?                      �?      �?                      �?�������?�������?      �?      �?              �?      �?              �?      �?              �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?              �?2'�����?3����?#��Q��?�(W��?j�V���?ˠT�x?�?|��|�?|���?�i��F�?GX�i���?      �?        �m۶m��?�$I�$I�?t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?              �?      �?      �?333333�?�������?              �?      �?                      �?(������?^Cy�5�?�������?�������?              �?      �?      �?۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?      �?        ��y��y�?�a�a�?      �?              �?      �?              �?      �?        ە�]���?�ڕ�]��?              �?UUUUUU�?UUUUUU�?      �?        333333�?ffffff�?              �?333333�?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?F]t�E�?�.�袋�?UUUUUU�?�������?              �?      �?                      �?�������?��U����?�\y@���?Ũ�oS��?�8�1�s�?�Ź�Q�?qG�wĭ?�;⎸#�?�������?�������?8��18�?�����?      �?        ;�;��?�؉�؉�?|���?|���?�?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?              �?h/�����?Lh/����?      �?        �;�;�?'vb'vb�?r�q��?�q�q�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?        �?<<<<<<�?�q�q�?9��8���?      �?      �?              �?      �?              �?                      �?]t�E�?t�E]t�?��y��y�?1�0��?(������?l(�����?      �?      �?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?              �?              �?              �?                      �?(�����?���k(�?      �?                      �?�B!��?���{��?h/�����?���Kh�?      �?      �?�q�q�?��8��8�?F]t�E�?]t�E�?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?                      �?              �?              �?              �?      �?      �?F]t�E�?/�袋.�?�q�q�?�q�q�?      �?                      �?      �?      �?              �?      �?        �������?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��-hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�Mh�h)h,K ��h.��R�(KM��h��B�C         p                    �?�ܲ�}��?�           ��@               M                    �?R�|[��?�            `w@              $                    �?�׺W4�?�            Pr@                                  �?���\=y�?�             k@                                 �c@      �?z             h@                                  �O@0G���ջ?D             Z@                                  @M@�x�E~�?;            @V@                                  �G@�}��L�?2            �R@        	       
                   �b@Pa�	�?            �@@       ������������������������       �                     =@                                   �?      �?             @        ������������������������       �                      @                                  o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@                                   ^@@4և���?	             ,@        ������������������������       �                     "@                                   �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  @t@������?	             .@                               ����?r�q��?             (@                                   `Q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@                                  Pc@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        6             V@                #                    l@�q�����?             9@        !       "                   pb@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     &@        %       4                    �K@���=A�?-             S@       &       /                   �?��k=.��?            �G@       '       .                   i@�L���?            �B@        (       -                    �?���!pc�?             &@       )       ,                    �?�����H�?             "@       *       +                   `^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@        0       3                 ����?���Q��?             $@       1       2                   @]@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        5       6                    @L@П[;U��?             =@        ������������������������       �                     @        7       B                    �?�q�����?             9@        8       9                   �`@�q�q�?             (@        ������������������������       �                      @        :       ;                   �c@�z�G��?             $@        ������������������������       �                     @        <       =                   �_@      �?             @        ������������������������       �                      @        >       A                    �?      �?             @       ?       @                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        C       F                    �?�n_Y�K�?             *@        D       E                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        G       H                    ]@���|���?             &@        ������������������������       �                      @        I       L                   �b@�<ݚ�?             "@       J       K                    U@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        N       e                   �b@������?6            @T@       O       `                    �?     8�?(             P@        P       _       	             �?�G�z��?             4@       Q       R                 ����?ҳ�wY;�?             1@        ������������������������       �                     @        S       ^                    �?d}h���?             ,@       T       [                    �?8�Z$���?             *@       U       V                    �?ףp=
�?             $@        ������������������������       �                      @        W       Z                    �?      �?              @        X       Y                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        \       ]                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        a       d                    U@���7�?             F@        b       c                   �`@      �?	             0@       ������������������������       �                     ,@        ������������������������       �                      @        ������������������������       �                     <@        f       o       	             �?j���� �?             1@       g       j                   �o@      �?             ,@        h       i                    �H@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        k       l                    �?�q�q�?             "@        ������������������������       �                      @        m       n                   pf@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        q       �                    �F@��A���?�            �v@        r       �                    �?���3�E�?&             J@        s       ~                 ����?      �?             8@        t       }                    �?�<ݚ�?             "@       u       x                   �`@      �?              @        v       w                   ``@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        y       z                    �D@r�q��?             @       ������������������������       �                     @        {       |       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               �                    �?�q�q�?
             .@       �       �       	             �?����X�?	             ,@       �       �                   �v@"pc�
�?             &@       �       �                    �?ףp=
�?             $@        ������������������������       �                      @        �       �       
             �?      �?              @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �? �Cc}�?             <@       �       �                   pb@�>����?             ;@       ������������������������       �                     3@        �       �                   �b@      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        �       �                    @C@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   a@��2(&�?�            @s@       �       �       
             �?���N8�?�            @j@       �       �                   `[@�]0��<�?w            �f@        ������������������������       �        &            �J@        �       �                    @Q@P�2E��?Q            @`@       �       �                 pff�?�m(']�?O            �_@        �       �                   P`@�C��2(�?            �@@       �       �                    �? 	��p�?             =@       �       �                   �[@ ��WV�?             :@        �       �                    �?؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             3@        �       �                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?`Ql�R�?<            �W@       �       �                    t@����e��?(            �P@       ������������������������       �        $             O@        �       �                    �?      �?             @       �       �                   �v@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?h�����?             <@       �       �                   �p@�}�+r��?             3@       �       �                   �n@ףp=
�?             $@       ������������������������       �                      @        �       �                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     "@        �       �                    �Q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?PN��T'�?             ;@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�8��8��?             8@       �       �                   p`@���N8�?             5@        �       �                     N@�����H�?             "@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             (@        �       �                   Pb@�q�q�?             @        ������������������������       �                     �?        �       �                 hff @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�J��%�?B            �X@       �       �                   �?�q���?"             H@        �       �                    `@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �q@�q�q�?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��
ц��?            �C@       �       �                    �M@|��?���?             ;@       �       �                    �?p�ݯ��?             3@       �       �       
             �?��S���?             .@        �       �                   Pd@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ����?�<ݚ�?             "@        ������������������������       �                     @        �       �                   �a@���Q��?             @        ������������������������       �                     �?        �       �                   pb@      �?             @        ������������������������       �                     �?        �       �                   @c@�q�q�?             @        ������������������������       �                     �?        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   `]@�q�q�?	             (@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                    d@����X�?             @       �       �                   0n@r�q��?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                         �c@j�q����?              I@       �                         �a@�Ra����?             F@        �                          �?�<ݚ�?             2@                               ����?և���X�?             @                                �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@                              hff�? ��WV�?             :@                                `g@z�G�z�?             @        ������������������������       �                     @        	      
                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@                                 �N@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �t�b�A#     h�h)h,K ��h.��R�(KMKK��hi�B�  ����u��?/�E��?0G��/�?�q��+��?:f���M�?gB����?�a��zX�?��Tx*<�?      �?      �?vb'vb'�?�؉�؉�?����G�?p�\��?�_,�Œ�?O贁N�?|���?|���?      �?              �?      �?      �?              �?      �?              �?      �?              �?        n۶m۶�?�$I�$I�?      �?        �������?�������?      �?                      �?wwwwww�?�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �p=
ף�?���Q��?�$I�$I�?۶m۶m�?              �?      �?              �?        ��P^Cy�?�P^Cy�?g���Q��?br1���?}���g�?L�Ϻ��?F]t�E�?t�E]t�?�q�q�?�q�q�?�������?UUUUUU�?              �?      �?              �?                      �?      �?        �������?333333�?�$I�$I�?۶m۶m�?      �?                      �?      �?        ��=���?�{a���?              �?�p=
ף�?���Q��?�������?�������?      �?        333333�?ffffff�?              �?      �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?ى�؉��?      �?      �?              �?      �?        ]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?      �?              �?      �?                      �?{	�%���?B{	�%��?      �?     ��?�������?�������?�������?�������?      �?        ۶m۶m�?I�$I�$�?;�;��?;�;��?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        F]t�E�?�.�袋�?      �?      �?              �?      �?                      �?�������?ZZZZZZ�?      �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        DDDDDD�?�������?b'vb'v�?O��N���?      �?      �?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?%I�$I��?h/�����?�Kh/��?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        t�E]t�?��.���?�a�a�?��y��y�?;ڼOqɠ?\2�h��?              �?z�z��?_�^��?
�B�P(�?����z��?F]t�E�?]t�E�?�{a���?������?;�;��?O��N���?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        W�+�ɕ?}g���Q�?|���?�>����?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?�m۶m��?(�����?�5��P�?�������?�������?              �?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?h/�����?&���^B�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�a�a�?��y��y�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?9/����?c}h���?�������?�������?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?�;�;�?�؉�؉�?{	�%���?	�%����?Cy�5��?^Cy�5�?�������?�?�������?UUUUUU�?      �?                      �?�q�q�?9��8���?              �?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?�������?�������?      �?              �?      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        
ףp=
�?=
ףp=�?]t�E�?]t�E]�?�q�q�?9��8���?�$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?                      �?;�;��?O��N���?�������?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�;GhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��B�;         �       	             �?znt��s�?�           ��@              �                    �?*|�� �?t           ��@              b                 ����?P�%f��?S           ��@               E                    �?~|z����?�            �p@              &                    @K@6��f�?`            @c@                                  �?�j�@�?:            �W@        ������������������������       �                     @@               #                     H@��s����?&            �O@       	                           �?>��C��?            �E@        
                          0n@��2(&�?             6@       ������������������������       �        
             0@                                  @c@      �?             @        ������������������������       �                     @        ������������������������       �                     @                                  �X@�q�q�?             5@        ������������������������       �                     �?                                   �?�z�G��?             4@                                   �?X�<ݚ�?             "@                                  `\@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   ^@z�G�z�?             @                                 �^@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?               "                 433�?"pc�
�?             &@              !                    �?ףp=
�?             $@                                   @D@؇���X�?             @                                  �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        $       %                    �?ףp=
�?
             4@       ������������������������       �        	             2@        ������������������������       �                      @        '       (                    �L
�q��?&            �M@        ������������������������       �                     @        )       B                   `c@Dc}h��?%             L@       *       =                    �?�<ݚ�?            �F@       +       6       
             �?�ݜ�?            �C@       ,       5                    �?�S����?             3@       -       4                    �?z�G�z�?             .@       .       1                   �d@؇���X�?             ,@       /       0                    U@�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        2       3                   f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        7       8                   `a@ףp=
�?             4@       ������������������������       �                     ,@        9       <                    �?�q�q�?             @        :       ;                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        >       A                    �?r�q��?             @        ?       @                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        C       D                    �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        F       W                    �?�MI8d�?B            �[@       G       P                 ����?��|���?4             V@       H       O                    �?`2U0*��?+            �R@       I       N                    @E@ "��u�?             I@        J       M                    �?�θ�?             *@        K       L                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                    �B@        ������������������������       �                     9@        Q       R                    X@�θ�?	             *@        ������������������������       �                      @        S       V                   `_@�C��2(�?             &@        T       U                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        X       Y                    �?��<b���?             7@        ������������������������       �                     @        Z       a                    �?�}�+r��?             3@       [       `                    �?@4և���?             ,@       \       ]       
             �?      �?              @       ������������������������       �                     @        ^       _                   Pm@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        c       �                    �?��%�V��?�            0q@        d       �                 ��� @�n_Y�K�?)            @P@       e       t                    �?�q���?              H@        f       m       
             �?�q�q�?             8@        g       h                    �?�q�q�?             @        ������������������������       �                     @        i       j                    �?�q�q�?             @        ������������������������       �                     �?        k       l                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        n       q                 033�?r�q��?             2@       o       p                   �Z@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        r       s                     H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        u       v                    �?�q�q�?             8@        ������������������������       �                     @        w       ~                    �?�����H�?             2@       x       }                    �M@��S�ۿ?             .@        y       |                    �?z�G�z�?             @       z       {                   Xq@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@               �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             1@        �       �                    �?ףp=
�?�            @j@       �       �                    �?�9��~�?_            �a@        �       �                    �?�Z��L��?.            �Q@        �       �                   xu@�E��ӭ�?             2@       ������������������������       �                     (@        �       �                    b@r�q��?             @        ������������������������       �                     @        �       �                    @O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �? �h�7W�?#            �J@       �       �                   Pr@ �q�q�?             H@       �       �                 033@ ���J��?            �C@       ������������������������       �                     ?@        �       �                   pk@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �r@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ����?z�G�z�?             @        �       �                    c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@�ӭ�a��?1             R@       �       �                    @H@���*�?*             N@        �       �                    �G@���|���?	             &@       ������������������������       �                     @        �       �                   �]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �a@؇���X�?!            �H@       �       �                    g@z�G�z�?             D@        �       �                   �^@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �b@     ��?             @@       ������������������������       �                     9@        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                    �K@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     (@        �       �                    �?0�,���?)            �P@       ������������������������       �        $            �L@        �       �                    Z@z�G�z�?             $@        �       �                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �C@���c���?!             J@        ������������������������       �                     �?        �       �                   �U@�t����?             �I@        ������������������������       �                     �?        �       �                    �?ףp=
�?             I@       �       �                    �?Du9iH��?            �E@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                    �L@z�G�z�?             @        ������������������������       �                     @        �       �                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   8r@г�wY;�?             A@       ������������������������       �                     >@        �       �                    �?      �?             @       �       �                    �R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?����X�?             @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @L@�Z��L��?_            �a@       �       �                   �g@ 7���B�?J             [@       �       �                    �? 5x ��?I            �Z@       �       �                    �?�ջ����?F             Z@       ������������������������       �        >            @W@        �       �                    @I@�C��2(�?             &@        ������������������������       �                     @        �       �                    �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @F@�q�q�?             @        ������������������������       �                     �?        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ҳ�wY;�?             A@       �       �                    _@�+$�jP�?             ;@        �       �                     Q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �u@���}<S�?             7@       �       �                    @M@���7�?             6@        �       �                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             1@        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ����?��}t��?���g��?��L��?�`�`�?�O��O��?�	�[���?��sHM0�?g�'�Y�?�cj`��?T��8��?�a�+�?      �?        z��y���?�a�a�?$�;��?qG�w��?��.���?t�E]t�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?ffffff�?333333�?r�q��?�q�q�?      �?      �?              �?      �?        �������?�������?      �?      �?      �?                      �?      �?        /�袋.�?F]t�E�?�������?�������?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?                      �?�������?�������?      �?                      �?��V'�?�pR���?              �?�$I�$I�?۶m۶m�?9��8���?�q�q�?\��[���?�i�i�?(������?^Cy�5�?�������?�������?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?F]t�E�?]t�E]�?              �?      �?        L�Ϻ��?��L���?颋.���?F]t�E�?{�G�z�?���Q��?���Q��?�G�z�?�؉�؉�?ى�؉��?      �?      �?              �?      �?                      �?              �?              �?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?      �?      �?              �?      �?              �?        ��Moz��?��,d!�?      �?        (�����?�5��P�?�$I�$I�?n۶m۶�?      �?      �?              �?      �?      �?              �?      �?                      �?              �?i�V1i�?�:[����?ى�؉��?;�;��?�������?�������?�������?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�������?UUUUUU�?�������?�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?�?�������?�������?�������?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?�U0K��?��3m���?��Vؼ?���.�d�?r�q��?�q�q�?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?"5�x+��?��sHM0�?UUUUUU�?�������?�A�A�?��-��-�?              �?      �?      �?      �?                      �?�q�q�?�q�q�?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?�8��8��?�q�q�?wwwwww�?""""""�?F]t�E�?]t�E]�?              �?�������?�������?              �?      �?        �$I�$I�?۶m۶m�?ffffff�?ffffff�?      �?      �?              �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?                      �?              �?g��1��?Ez�rv�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�;�;�?;�;��?      �?        �?<<<<<<�?      �?        �������?�������?w�qGܱ?qG�w��?�q�q�?9��8���?      �?              �?      �?�������?�������?              �?      �?      �?              �?      �?                      �?�?�?              �?      �?      �?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?���.�d�?��Vؼ?	�%����?h/�����?7��XQ�?�@�Ե�?;�;��?;�;��?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�������?�������?/�����?B{	�%��?      �?      �?              �?      �?        ӛ���7�?d!Y�B�?�.�袋�?F]t�E�?�������?�������?              �?      �?              �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�a{8hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK�h��B�<         b                   P`@�_y���?�           ��@               O       	             �?\�f<t�?�            @t@              6                   �a@���7��?�             r@              #                    �?>���$��?            �g@                               pff�?��S�ۿ?h            �b@                                  �_@(2��R�?,            �M@        ������������������������       �                     =@               	                 ����?������?             >@        ������������������������       �                     @        
                           �K@�LQ�1	�?             7@        ������������������������       �                     @                                  �`@��.k���?             1@                                    P@�<ݚ�?             "@                                  �?      �?              @                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   �?      �?              @       ������������������������       �                     @                                  �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                    �Q@p�C��?<            �V@                                  �J@�|���?:             V@                                   @J@ �q�q�?             8@       ������������������������       �                     6@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        *             P@        !       "                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        $       5                 033�?R���Q�?             D@       %       (                    U@4?,R��?             B@        &       '                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        )       *                   �X@     ��?             @@        ������������������������       �                     �?        +       .                    �E@`Jj��?             ?@        ,       -                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        /       4                    W@h�����?             <@        0       3                   @\@r�q��?             @       1       2                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                     @        7       J       
             �?ףp=
�?E             Y@       8       I                    �R@����?:            �U@       9       B                    �?�IєX�?9            @U@       :       ?                   0`@ ���J��?3            �S@       ;       >                    �?`׀�:M�?0            �R@        <       =                   pb@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        ,            @Q@        @       A                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        C       D                    �?և���X�?             @        ������������������������       �                     �?        E       H                   �c@�q�q�?             @       F       G                   �\@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        K       N                    �M@�θ�?             *@       L       M                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        P       W                   �?��.k���?             A@       Q       R                   �b@��S�ۿ?
             .@       ������������������������       �                     (@        S       V                    �?�q�q�?             @       T       U                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        X       a                    �?���y4F�?             3@       Y       \                    �?      �?             0@        Z       [                   `c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ]       `                    �?�8��8��?             (@        ^       _                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        c       �                    @L@l�C�o��?           �y@       d       m                   �^@      �?�             q@        e       l       	             �?�㙢�c�?             7@       f       k                   �a@��2(&�?             6@        g       h                    �?�q�q�?             "@        ������������������������       �                     �?        i       j                   �a@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     �?        n       �                    �?�>��_;�?�             o@       o       �                   �{@��UV�?�            �j@       p       �                    �?�����?�            `j@       q       |                    �?h�|�6�?g            @e@        r       s                    �?���C��?"            �J@        ������������������������       �                     6@        t       y                    �?�n`���?             ?@       u       v                   `q@�nkK�?             7@       ������������������������       �                     5@        w       x                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        z       {                     G@      �?              @        ������������������������       �                     @        ������������������������       �                     @        }       ~                    �?�6H�Z�?E            @]@       ������������������������       �        4            �V@               �                    �? ��WV�?             :@        ������������������������       �                     @        �       �                   �d@���N8�?             5@       ������������������������       �        	             0@        �       �                    �G@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�>$�*��?            �D@       �       �                 ����?:ɨ��?            �@@       �       �                   �d@V�a�� �?             =@       �       �                    �?ҳ�wY;�?             1@       �       �       	             �?d}h���?             ,@        �       �                   d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     C@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �        	             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?b�2�tk�?             B@       �       �                   �l@���!pc�?             6@       �       �                    �?�eP*L��?	             &@        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �J@����X�?             @       �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �c@և���X�?             ,@        ������������������������       �                     @        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �       
             �?z�G�z�?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �Z@�û��|�?X            @a@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �`@z���ȋ�?T            @`@        �       �                 ��� @��+7��?              G@       �       �                    �?�q�q�?             B@       �       �                 ����?X�<ݚ�?             ;@        �       �                    �M@�eP*L��?	             &@        �       �                 ����?z�G�z�?             @        ������������������������       �                      @        �       �                     M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   (r@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   `m@      �?
             0@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     "@        ������������������������       �                     $@        �       �                    �?�q�q�?4             U@       �       �                 ����? s�n_Y�?             J@       �       �                    �M@\X��t�?             7@        �       �                    �?      �?              @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ����?��S���?             .@        ������������������������       �                      @        �       �                 ����?�n_Y�K�?
             *@        ������������������������       �                      @        �       �                   `a@�eP*L��?             &@        ������������������������       �                     �?        �       �                    �O@���Q��?             $@       �       �                   @e@�q�q�?             "@       �       �                   `c@և���X�?             @       �       �                   �p@�q�q�?             @        ������������������������       �                      @        �       �                   �u@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    c@XB���?             =@       ������������������������       �        
             3@        �       �                 `ff@ףp=
�?             $@        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@      �?             @@        �       �                    �?@4և���?             ,@       �       �                    �?ףp=
�?	             $@       ������������������������       �                     @        �       �                 ��� @      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   pd@b�2�tk�?             2@        �       �                   `r@�<ݚ�?             "@       �       �                   d@�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  V�.�#��?աh6n��?&���^B�?��Kh/�?_*h����?h���V_�?�%N���?��v�@�?�?�������?'u_[�?=�"h8��?              �?�?wwwwww�?              �?d!Y�B�?Nozӛ��?              �?�?�������?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?        h�h��?��K��K�?F]t�E�?��.���?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�8��8��?r�q��?      �?      �?      �?                      �?      �?      �?              �?���{��?�B!��?UUUUUU�?UUUUUU�?      �?                      �?�m۶m��?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?�������?�������?/�I���?��֡�l�?�?�?�A�A�?��-��-�?к����?��L��?�������?�������?              �?      �?                      �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �؉�؉�?ى�؉��?      �?      �?              �?      �?                      �?�������?�?�������?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        (������?6��P^C�?      �?      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?#t/B�"�?��{��?      �?      �?d!Y�B�?�7��Mo�?t�E]t�?��.���?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        &sp��?h3�?R0�?2~�ԓ��?6��9�?��^Fb5�?`�
��T�?�������?�?\�琚`�?"5�x+��?      �?        �9�s��?�c�1��?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        �������?���?      �?        O��N���?;�;��?      �?        ��y��y�?�a�a�?      �?        �������?�������?      �?                      �?�18���?�����?N6�d�M�?e�M6�d�?��{a�?a���{�?�������?�������?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?]t�E�?F]t�E�?              �?      �?                      �?      �?                      �?              �?              �?9��8���?�8��8��?t�E]t�?F]t�E�?t�E]t�?]t�E�?      �?      �?              �?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?              �?�q�q�?�q�q�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��,d!�?8��Moz�?      �?      �?      �?                      �?7r#7r#�?�Fn�Fn�?Y�B��?zӛ����?UUUUUU�?UUUUUU�?�q�q�?r�q��?t�E]t�?]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?              �?�������?�������?;�;��?�;�;�?��Moz��?!Y�B�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�������?              �?;�;��?ى�؉��?      �?        t�E]t�?]t�E�?              �?333333�?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?                      �?�{a���?GX�i���?              �?�������?�������?      �?      �?              �?      �?                      �?      �?      �?n۶m۶�?�$I�$I�?�������?�������?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        �8��8��?9��8���?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ ��#hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKυ�h��B�3         |                    �?"�\�&U�?�           ��@              A                    �?Z�0���?           pz@               (       
             �?���<��?l            �e@                                  �?     8�?O             `@                                `ff�?�q�q�?	             (@        ������������������������       �                      @                                  @_@z�G�z�?             $@        ������������������������       �                     @        	       
                   �T@      �?             @        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                833�?Riv����?F             ]@        ������������������������       �                    �G@                                  �^@��+7��?*            @Q@        ������������������������       �                     9@               #                    �?8�A�0��?             F@              "                   �a@��Zy�?            �C@                                  @I@�f7�z�?             =@                                  @f@�q�q�?             (@                     	             �?���!pc�?             &@       ������������������������       �                     @                                  Po@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?������?             1@        ������������������������       �                      @                                   `@X�<ݚ�?             "@        ������������������������       �                     @                !                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        $       %                    �?z�G�z�?             @        ������������������������       �                      @        &       '                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        )       *                 ����?z�J��?            �G@        ������������������������       �                      @        +       6                 `ff�?�n_Y�K�?            �C@       ,       1                    m@�㙢�c�?             7@       -       0                    �H@      �?	             0@        .       /                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        2       5                     P@և���X�?             @       3       4                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        7       8                    �?     ��?             0@        ������������������������       �                      @        9       >                   �c@d}h���?
             ,@       :       =                     H@�����H�?             "@        ;       <                    m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ?       @                   �_@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        B       u                    �?X��Oԣ�?�             o@       C       t                   h@$Nz�{�?�             k@       D       c                   �?�>����?�             k@       E       T                    �?���r�?x             f@       F       I                   `^@ ��ʻ��?\             a@        G       H                    ^@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        J       K                   `a@��d��?O             ^@       ������������������������       �        =            �W@        L       S                   �a@`2U0*��?             9@        M       N                    �?��S�ۿ?	             .@        ������������������������       �                      @        O       P                    �?$�q-�?             *@        ������������������������       �                     �?        Q       R                   xt@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �        	             $@        U       \                    �?,���i�?            �D@       V       [                   �i@�IєX�?             A@        W       X                    �?r�q��?             (@        ������������������������       �                      @        Y       Z                   @h@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        ]       ^                    �?և���X�?             @        ������������������������       �                      @        _       `                   g@���Q��?             @        ������������������������       �                      @        a       b                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        d       s                    �?�θ�?            �C@       e       p                   �_@¦	^_�?             ?@        f       g                    �?�n_Y�K�?             *@        ������������������������       �                      @        h       o       
             �?�eP*L��?	             &@       i       l       	             �?�q�q�?             "@       j       k                 ����?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        m       n                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        q       r                 ���@�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        v       {                     P@f���M�?             ?@       w       x                    �?�θ�?             :@       ������������������������       �                     3@        y       z                    `@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        }       �                    �?�q�޴�?�            ps@        ~       �                   `c@��
ц��?            �C@              �                    �?      �?             A@        ������������������������       �                     "@        �       �                    �J@`�Q��?             9@        �       �                    �?��
ц��?             *@        ������������������������       �                      @        �       �                    Z@���|���?             &@        ������������������������       �                      @        �       �                   �`@�<ݚ�?             "@       �       �                 ����?�q�q�?             @       �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    \@�8��8��?             (@        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ����?���� �?�             q@        �       �                    �?      �?(             Q@        �       �                   `d@`՟�G��?             ?@       �       �                   `a@��+7��?             7@       �       �                    �?      �?
             0@       �       �                     L@      �?             (@        ������������������������       �                     @        �       �                   �Z@      �?              @       �       �                   �a@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �L@�L���?            �B@        ������������������������       �        	             1@        �       �                    @M@R���Q�?             4@        �       �                   �l@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?��S�ۿ?
             .@       �       �                 ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���'Z��?�            �i@       �       �                   �`@P���Q�?�             i@       �       �                   @s@`#`��k�?b             c@       ������������������������       �        W            `a@        �       �                    �?؇���X�?             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?
             *@        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���	@t/*�?            �G@       �       �                   �Z@� ��1�?            �D@        ������������������������       �                     @        �       �                   �^@�?�'�@�?             C@        �       �                   �\@�q�q�?             (@        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @M@ ��WV�?             :@       ������������������������       �                     .@        �       �                    �M@�C��2(�?             &@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                 ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��j��`�?:�J;�O�?�b[ox�?�:I!��?��Ħ��?�����?      �?     ��?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?	�=����?>�����?              �?Y�B��?zӛ����?              �?/�袋.�?颋.���?\��[���?� � �?O#,�4��?a���{�?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?      �?        xxxxxx�?�?      �?        r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?AL� &W�?}g���Q�?              �?;�;��?ى�؉��?�7��Mo�?d!Y�B�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?              �?      �?      �?        ۶m۶m�?I�$I�$�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?�������?333333�?              �?      �?        c�1�c�?�s�9�?��u�:~�?�8P(�?�Kh/��?h/�����?�
���?�^o�?�?�������?�?      �?      �?      �?                      �?�������?�?      �?        ���Q��?{�G�z�?�������?�?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �����?8��18�?�?�?�������?UUUUUU�?      �?        �������?�������?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?ى�؉��?�؉�؉�?��Zk���?�RJ)���?ى�؉��?;�;��?              �?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ��8��8�?�q�q�?      �?                      �?      �?                      �?��RJ)��?��Zk���?ى�؉��?�؉�؉�?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?�g��p��?f�Σ�?�؉�؉�?�;�;�?      �?      �?      �?        {�G�z�?��(\���?�;�;�?�؉�؉�?              �?]t�E]�?F]t�E�?              �?9��8���?�q�q�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?�������?�������?              �?      �?        <<<<<<�?xxxxxx�?      �?      �?�s�9��?�1�c��?Y�B��?zӛ����?      �?      �?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?        L�Ϻ��?}���g�?              �?333333�?333333�?�������?333333�?              �?      �?        �?�������?      �?      �?              �?      �?                      �?PPPPPP�?�������?�������?ffffff�?p�pŊ?@�?��?              �?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?�������?      �?                      �?W�+���?�;����?������?������?      �?        y�5���?������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?;�;��?O��N���?              �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�?�hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��B@6         `                    �?�#i����?�           ��@               A                    �?Te�$��?�             u@               0                   �c@P����?J            �\@              #                   pb@�~�4_��?8             V@                                  �?д>��C�?(             M@                                  @_@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        	                           �?^�!~X�?$            �J@        
                        033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     @               "                    �?�r����?            �F@              !                   (s@"pc�
�?            �@@                                 `@     ��?             @@       ������������������������       �                     1@                                    �?�q�q�?             .@                                 �a@      �?	             $@                                   �?      �?             @                                   C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                      
             �?�q�q�?             @        ������������������������       �                      @                                  �b@      �?             @        ������������������������       �                     �?                                  �\@�q�q�?             @        ������������������������       �                     �?                                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        $       '                    ]@�z�G��?             >@        %       &                     P@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        (       -                    �?z�G�z�?             9@       )       *                    �M@�����H�?	             2@       ������������������������       �                     &@        +       ,       
             �?����X�?             @        ������������������������       �                     @        ������������������������       �                      @        .       /                     Q@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        1       :                    @�θ�?             :@       2       7                    �?"pc�
�?             6@       3       4                   @a@�KM�]�?             3@       ������������������������       �        
             0@        5       6                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        8       9                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ;       @                    �?      �?             @       <       ?                   �e@�q�q�?             @       =       >                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        B       M                    �? �Cc��?�             l@        C       J                     R@f>�cQ�?(            �N@       D       E                    �?�KM�]�?&            �L@        ������������������������       �                     3@        F       I                   �c@�S����?             C@       G       H                 hff@�����H�?             B@       ������������������������       �                     @@        ������������������������       �                     @        ������������������������       �                      @        K       L                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        N       _                    �?������?e            `d@       O       T                   @[@�g<a�?`            @c@        P       S                    c@؇���X�?             @        Q       R                   �_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        U       ^                   �c@@�E�x�?Y            `b@       V       W                    @L@P��BNֱ?3            �T@       ������������������������       �        &             O@        X       ]                   �s@؇���X�?             5@       Y       \                   �_@ףp=
�?             4@        Z       [                   �p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             0@        ������������������������       �                     �?        ������������������������       �        &             P@        ������������������������       �                     "@        a       �                    �?*S%��?�            �x@       b       �                    �M@4V��X�?�            `q@       c       p                   `\@�Lt�?w            �f@        d       m                    �?     ��?             @@       e       f                   �i@p�ݯ��?             3@        ������������������������       �                     @        g       l                 033@�q�q�?             (@       h       k                   �m@X�<ݚ�?             "@        i       j                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        n       o                    q@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        q       �                    �?.�W����?a            �b@        r       s                   �]@���|���?!            �K@        ������������������������       �                     @        t       �                    b@θ	j*�?             J@       u       ~                   �g@��Q���?             D@        v       w                    �?X�<ݚ�?             2@        ������������������������       �                      @        x       y                     G@z�G�z�?             $@        ������������������������       �                     �?        z       }                   @E@�����H�?             "@        {       |                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               �                    �G@���7�?             6@        �       �                   �k@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                    �?      �?             (@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�"�q��?@            �W@       �       �                    _@�o��gn�?8            �T@        �       �                     H@�z�G��?             4@        ������������������������       �                     @        �       �                   �o@���Q��?             .@       ������������������������       �                      @        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�[|x��?-            �O@        �       �                    �J@      �?              @       �       �                    �I@���Q��?             @       �       �                 ����?      �?             @        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�1�`jg�?%            �K@       �       �                    �? �q�q�?             H@       �       �                   �a@�IєX�?             A@       �       �                    @M@�KM�]�?             3@       ������������������������       �                     .@        �       �                   b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             .@        ������������������������       �                     ,@        �       �                   �Y@؇���X�?             @        ������������������������       �                     @        �       �                   `c@�q�q�?             @       �       �                   @\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    c@      �?             (@       �       �                   �`@      �?              @        ������������������������       �                      @        �       �                   �k@�q�q�?             @        ������������������������       �                     �?        �       �                   pf@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �V@     ��?6             X@        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    l@xP�Fֺ�?2            @V@        �       �                    �?��<b���?             G@        �       �                    �?      �?
             0@       �       �                 @33�?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     >@        �       �                 ����? qP��B�?            �E@        �       �                    ^@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �A@        �       �                   Pz@����˵�?I            �]@       �       �                    �I@ T���v�?G            @\@        �       �                    �?ȵHPS!�?             :@        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�}�+r��?             3@       ������������������������       �        	             *@        �       �                   �_@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        6            �U@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �t�b�@     h�h)h,K ��h.��R�(KK�KK��hi�B�  �5�;���?%e��?d���+��?8�Z$���?Q^Cy��?�P^Cy�?��.���?]t�E�?|a���?a���{�?333333�?�������?      �?                      �?�	�[���?�}�	��?      �?      �?      �?                      �?�?�������?F]t�E�?/�袋.�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?                      �?333333�?ffffff�?�������?�������?              �?      �?        �������?�������?�q�q�?�q�q�?              �?�$I�$I�?�m۶m��?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ى�؉��?�؉�؉�?/�袋.�?F]t�E�?�k(���?(�����?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?I�$I�$�?n۶m۶�?��!XG�?�u�y���?�k(���?(�����?      �?        (������?^Cy�5�?�q�q�?�q�q�?      �?                      �?              �?      �?      �?              �?      �?        �x�%�6�?)��I� �?���8+�?�cj`?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        և���X�?9/���?��FS���?���ˊ��?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?              �?        �v�ļ�?;Cb�ΐ�?���n��?'!����?y��x���?D8�C8��?      �?      �?Cy�5��?^Cy�5�?              �?�������?�������?�q�q�?r�q��?�������?�������?      �?                      �?              �?      �?        �؉�؉�?;�;��?      �?                      �?0��b�/�?贁N��?]t�E]�?F]t�E�?              �?�؉�؉�?�N��N��?333333�?�������?�q�q�?r�q��?              �?�������?�������?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �.�袋�?F]t�E�?      �?      �?      �?      �?              �?      �?              �?              �?              �?      �?              �?      �?      �?              �?      �?        |n�S���?a�+F�?�7�:���?rY1P��?333333�?ffffff�?              �?�������?333333�?              �?۶m۶m�?�$I�$I�?      �?                      �?EQEQ�?]�u]�u�?      �?      �?�������?333333�?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?�־a�?A��)A�?UUUUUU�?�������?�?�?(�����?�k(���?              �?      �?      �?              �?      �?                      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?              �?      �?�$I�$I�?۶m۶m�?      �?                      �?�я~���?�.p��?��Moz��?��,d!�?      �?      �?]t�E�?F]t�E�?              �?      �?                      �?              �?�}A_З?��}A�?      �?      �?      �?      �?      �?                      �?              �?              �?��/���?W'u_�?4��A�/�?6h�e�&�?�؉�؉�?��N��N�?�$I�$I�?�m۶m��?      �?                      �?(�����?�5��P�?              �?UUUUUU�?�������?      �?                      �?              �?333333�?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	Ͳ$hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�?         |                    @L@�$���?�           ��@              C                    �?RA��lZ�?           �y@               :                    �?�ُT�?            �h@                                 Pi@�k�'7��?i            `e@                      	             �?,�+�C�?$            �K@                                  �?`'�J�?!            �I@                                   �?z�G�z�?             $@       ������������������������       �                     @        	       
                   @Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �D@                                `ff�?      �?             @        ������������������������       �                      @        ������������������������       �                      @               /                   q@^l��[B�?E             ]@                                  _@<ݚ)�?+             R@                                  @c@�q�q�?             8@                                  �?��S���?             .@                                 �\@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                    D@�<ݚ�?             "@        ������������������������       �                     �?                                  e@      �?              @                                 Pl@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               &                 ����?r�q��?             H@                !                   pi@�����?             3@        ������������������������       �                      @        "       #                   l@������?
             1@        ������������������������       �                     $@        $       %                   �l@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        '       *                    �? 	��p�?             =@        (       )                     K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        +       ,       
             �? ��WV�?             :@       ������������������������       �                     7@        -       .                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        0       9                    f@�C��2(�?             F@       1       2                   xt@��Y��]�?            �D@       ������������������������       �                     =@        3       4                    �?�8��8��?             (@        ������������������������       �                     @        5       8                     J@      �?              @       6       7                    �H@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ;       >                   �g@��>4և�?             <@        <       =                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ?       B                   �b@���!pc�?             6@        @       A                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             .@        D       U                    �?�e/
�?�             k@       E       R                   �g@P-�T6��?_            �b@       F       Q                    @@�E�x�?]            `b@       G       H       
             �? �й���?\            @b@       ������������������������       �        9             W@        I       J                    �? 7���B�?#             K@        ������������������������       �                     1@        K       P                   c@@-�_ .�?            �B@        L       M                   0n@�����H�?             2@       ������������������������       �                     $@        N       O                   �]@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                     �?        S       T                    �D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        V       m                    `@�	j*D�?*            @P@       W       f                   @^@     ��?             @@       X       a                    �?�q�q�?             8@       Y       Z                    @D@���y4F�?             3@        ������������������������       �                      @        [       `                   �q@�t����?             1@       \       ]                    �?      �?
             0@       ������������������������       �                     *@        ^       _                   a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        b       e                    �H@z�G�z�?             @       c       d                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        g       h                    �F@      �?              @        ������������������������       �                     @        i       l                    �?�q�q�?             @       j       k                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        n       u                    �?6YE�t�?            �@@       o       t                    �? �q�q�?             8@       p       q                    �?���N8�?             5@        ������������������������       �                     @        r       s                    �D@�X�<ݺ?
             2@        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     @        v       w                   �^@X�<ݚ�?             "@        ������������������������       �                      @        x       {                    �J@����X�?             @       y       z                 ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        }       �                    �?�c�Α�?�            �s@        ~       �                    �?��
ц��?R            @`@              �                   �d@:PZ(8?�?0            @R@        �       �                    �?b�2�tk�?             2@       �       �                    �?���|���?             &@       �       �       	             �?�q�q�?             @       �       �                    `Q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Hp@x��}�?%            �K@       �       �                    �M@�8��8��?             B@        �       �                    �?d}h���?
             ,@       �       �                   �`@���!pc�?             &@       �       �                 ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        �       �       	             �?�\��N��?             3@       �       �       
             �?�q�q�?
             .@       �       �                    �?�θ�?             *@        ������������������������       �                     @        �       �                    �?�q�q�?             "@       �       �                   p`@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?F�t�K��?"            �L@        ������������������������       �                      @        �       �                    @N@�2����?             �K@       �       �                    �?�q�q�?             ;@        ������������������������       �                     @        �       �                    �?�G�z��?             4@       �       �                   �n@X�Cc�?             ,@       �       �                   �V@�	j*D�?             *@        ������������������������       �                      @        �       �                    �?"pc�
�?             &@       �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                     M@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        �       �                   �x@PN��T'�?p            �g@       �       �                    �?$G$n��?m             g@        �       �                    �?      �?-             R@        �       �                 pff�?���!pc�?             &@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �Z@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `\@��.��?'            �N@        ������������������������       �                     8@        �       �       
             �?����>�?            �B@       �       �                 pff�?d}h���?             <@       �       �                 ����?ҳ�wY;�?             1@       �       �                    �?8�Z$���?             *@        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @]@�C��2(�?             &@        ������������������������       �                     @        �       �                   �n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    �N@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@ (��?@            @\@       �       �                    �?�f�¦ζ?<            �Z@        �       �                    �?H%u��?             9@       �       �                   �`@�8��8��?             8@       �       �                    �?���7�?             6@       �       �                    �?�8��8��?             (@       �       �       
             �?ףp=
�?             $@        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                 `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��Y��]�?.            �T@       �       �                    �?h㱪��?            �K@       ������������������������       �                    �C@        �       �                 ����?      �?
             0@        �       �                   `X@      �?              @        ������������������������       �                     �?        �       �                   `b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        �       �                   �c@�q�q�?             @       �       �                 `ff�?      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  �E$�~V�?�����?C��RF�?z���Zs�?�n-;�?zWd�4q�?Lg1��t�?-����b�?��)A��?�}��7��?�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        ��=���?�=�����?�8��8��?��8��8�?�������?�������?�������?�?�������?�������?              �?      �?              �?        9��8���?�q�q�?              �?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?�������?^Cy�5�?Q^Cy��?      �?        �?xxxxxx�?              �?�$I�$I�?۶m۶m�?      �?                      �?�{a���?������?UUUUUU�?UUUUUU�?      �?                      �?;�;��?O��N���?              �?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E�?������?8��18�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?              �?      �?                      �?      �?        ۶m۶m�?I�$I�$�?UUUUUU�?�������?      �?                      �?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?                      �?      �?        _B{	�%�?	�%��о?���t}��?�`Q�(X�?և���X�?9/���?����Ǐ�?����?      �?        	�%����?h/�����?      �?        S�n0E�?к����?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?                      �?      �?      �?      �?                      �?vb'vb'�?;�;��?      �?      �?UUUUUU�?UUUUUU�?6��P^C�?(������?              �?<<<<<<�?�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?      �?              �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?'�l��&�?e�M6�d�?�������?UUUUUU�?��y��y�?�a�a�?      �?        ��8��8�?�q�q�?              �?      �?              �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?�{a���?5�rO#,�?�؉�؉�?�;�;�?�W�^�z�?�P�B�
�?9��8���?�8��8��?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?pX���o�?A��)A�?UUUUUU�?UUUUUU�?I�$I�$�?۶m۶m�?F]t�E�?t�E]t�?�������?333333�?      �?                      �?      �?              �?              �?        �5��P�?y�5���?UUUUUU�?UUUUUU�?�؉�؉�?ى�؉��?              �?UUUUUU�?UUUUUU�?      �?      �?              �?�������?333333�?              �?      �?              �?              �?              �?        :��,���?1��t��?      �?        � O	��?��7�}��?UUUUUU�?UUUUUU�?              �?�������?�������?%I�$I��?�m۶m��?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?              �?h/�����?&���^B�?���L�?к����?      �?      �?F]t�E�?t�E]t�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ������?�����?              �?���L�?�u�)�Y�?۶m۶m�?I�$I�$�?�������?�������?;�;��?;�;��?      �?      �?              �?      �?        F]t�E�?]t�E�?              �?      �?      �?      �?                      �?      �?                      �?�q�q�?r�q��?              �?�������?�������?      �?              �?      �?              �?      �?        x�!���?H���?�Ե��?��4>2��?���Q��?)\���(�?UUUUUU�?UUUUUU�?F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?              �?        ������?8��18�?��)A��?־a���?              �?      �?      �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�J�	hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKŅ�h��B@1         R                    �?6������?�           ��@                                   @K@�x�W�?�             w@                                  �?T�y���?�            `j@                                  �?@�K�҈?d            �d@       ������������������������       �        a             d@                      
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        	                          �b@p�v>��?             �G@       
                           P@@4և���?             <@                                   Z@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     8@                                ����?p�ݯ��?             3@                               `ffֿ��
ц��?
             *@        ������������������������       �                      @                                   ]@�eP*L��?	             &@        ������������������������       �                     @                                  �d@      �?              @        ������������������������       �                      @        ������������������������       �                     @                                   b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?               I       	             �?�Zi`���?c            �c@              *                    �?2?74e��?N            @_@               )                    �?p9W��S�?             C@              (                 ��� @      �?             B@              '                    �?"pc�
�?            �@@              "                    d@V�a�� �?             =@               !                   �b@�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @        #       $                    �?���Q��?             $@       ������������������������       �                     @        %       &                    �M@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        +       B                    �?�q�q�?3            �U@       ,       =                    �?4�.�A�?#            �O@       -       8                   0a@      �?             F@       .       3                 @33�?�+e�X�?             9@        /       0                    �?      �?             @        ������������������������       �                     �?        1       2                   �]@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        4       5                   �]@؇���X�?             5@        ������������������������       �                     &@        6       7                   �U@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        9       <                    �?�S����?	             3@       :       ;                    �?�����H�?             2@       ������������������������       �                     0@        ������������������������       �                      @        ������������������������       �                     �?        >       A                    �L@���y4F�?
             3@        ?       @                 @33�?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        C       D                    �?      �?             8@        ������������������������       �                      @        E       H                 ����?     ��?
             0@        F       G                   `\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        J       O                     R@     ��?             @@       K       L                   �?��S�ۿ?             >@       ������������������������       �                     :@        M       N                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        P       Q                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       �                   �c@f>�cQ�?�            �v@       T       �       	             �?<�jX��?�            �s@       U       V                    Z@��v�u�?�            `r@        ������������������������       �                    �G@        W       f                    �?� � J��?�            �n@        X       _                 ����?���!pc�?             6@       Y       ^                   �`@�8��8��?
             (@        Z       [                    �?z�G�z�?             @        ������������������������       �                      @        \       ]                    b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        `       c                    �?      �?             $@       a       b                 ���@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        d       e                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        g       �                   P`@4���|��?�             l@        h       i                   �h@��E�wx�?E            �[@        ������������������������       �                    �F@        j       �                    �?F.< ?�?)            �P@       k       |                    �?x��}�?$            �K@        l       {                   pp@������?             >@       m       z                    �?��.k���?
             1@       n       s                    �K@���Q��?	             .@        o       p                   @^@      �?             @        ������������������������       �                      @        q       r                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        t       u                   `@���!pc�?             &@        ������������������������       �                      @        v       y                    �?�����H�?             "@       w       x                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        }       �                    �?z�G�z�?             9@        ~       �                    @L@���Q��?             @              �                    �?�q�q�?             @       �       �                   m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?ףp=
�?             4@       �       �                    [@r�q��?
             (@        ������������������������       �                     �?        �       �                    `@�C��2(�?	             &@        �       �                   `_@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?���U�?K            �\@        �       �                   �d@���}<S�?             7@       �       �                    �?���7�?             6@       ������������������������       �        
             ,@        �       �                   �?      �?              @        �       �                   pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 033�?p�C��?;            �V@        �       �                    �?      �?              @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   pa@��'�`�?5            �T@       ������������������������       �        +             Q@        �       �                 ����?��S�ۿ?
             .@        �       �                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?���Q��?             4@       �       �                   @j@      �?	             (@        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��WV��?             J@       �       �                    �?և���X�?            �A@       �       �                   �n@ �o_��?             9@       �       �                    �?�IєX�?
             1@       ������������������������       �                     ,@        �       �       	             �?�q�q�?             @       �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@      �?              @        �       �                   d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    `@z�G�z�?             $@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �r@@�0�!��?             1@       ������������������������       �        	             ,@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  ��X�5�?��S�$e�?�7��Mo�?d!Y�B�?&�k]���?�&��2�?���|��?�����x?      �?              �?      �?              �?      �?        ڨ�l�w�?L� &W�?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?        Cy�5��?^Cy�5�?�؉�؉�?�;�;�?              �?t�E]t�?]t�E�?              �?      �?      �?              �?      �?        UUUUUU�?�������?              �?      �?        �5��(S�?b��x�Y�?y�&1��?D�l����?�k(����?l(�����?      �?      �?/�袋.�?F]t�E�?��{a�?a���{�?�k(���?(�����?      �?                      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?UUUUUU�?UUUUUU�?��i��i�?�,˲,��?      �?      �?���Q��?R���Q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?333333�?ffffff�?      �?                      �?(������?^Cy�5�?�q�q�?�q�q�?      �?                      �?              �?(������?6��P^C�?�q�q�?r�q��?      �?                      �?              �?      �?      �?              �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?�������?�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?�u�y���?��!XG�?�x�YF�?�0�T<��?e�J��?`��!�?              �?i}��ַ?S���.�?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?333333�?�������?      �?                      �?�������?333333�?      �?                      �?�h$��W�?�r����?���+c��?	ą��@�?              �?6�d�M6�?��&�l��?A��)A�?pX���o�?�?wwwwww�?�?�������?�������?333333�?      �?      �?      �?              �?      �?              �?      �?        t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?UUUUUU�?�������?      �?                      �?              �?      �?                      �?�������?�������?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        �������?�������?UUUUUU�?�������?      �?        F]t�E�?]t�E�?�������?�������?              �?      �?                      �?              �?              �?p�}��?	�#����?d!Y�B�?ӛ���7�?F]t�E�?�.�袋�?              �?      �?      �?      �?      �?              �?      �?                      �?      �?        h�h��?��K��K�?      �?      �?      �?      �?      �?                      �?              �?��k���?1P�M��?              �?�?�������?      �?      �?              �?      �?                      �?�������?333333�?      �?      �?      �?              �?      �?              �?      �?              �?      �?      �?                      �?��N��N�?��؉���?�$I�$I�?۶m۶m�?
ףp=
�?�Q����?�?�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?�������?333333�?              �?      �?                      �?�������?ZZZZZZ�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��qhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK녔h��B�:         �                    �?�+	G�?�           ��@              _                    �?����/��?w           �@              R                    �?�C���\�?�            0s@              #                    �?�r����?�            �p@              "                   �g@`h���?            �g@                                 �c@f�1�?~             g@                                 @[@ qP��B�?v            �e@               	                   0n@$�q-�?	             *@       ������������������������       �                     "@        
                           @I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�O4R���?m            �c@                                  I@�1���܋?e            @b@                                  0`@ףp=
�?             $@                                  �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        _             a@                                   �?8�Z$���?             *@        ������������������������       �                     @                                  0i@����X�?             @        ������������������������       �                     @                                  �b@      �?             @       ������������������������       �                      @        ������������������������       �                      @               !                    �P@8�Z$���?             *@                                  �?�8��8��?             (@       ������������������������       �                      @                                    @N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        $       I                 ����?�w���?1            @T@       %       B                   �q@���!pc�?&            �P@       &       =                   �l@j�q����?              I@       '       6                    �?      �?             @@       (       5                 @33�?H%u��?             9@       )       2                   �k@��2(&�?             6@       *       /                   �c@ףp=
�?             4@       +       ,                    �?      �?             0@       ������������������������       �        	             *@        -       .                     P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        0       1                   Pd@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        3       4                    @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        7       8                   g@����X�?             @        ������������������������       �                      @        9       <                    �?���Q��?             @       :       ;                   Pa@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        >       A                    `@�X�<ݺ?
             2@        ?       @                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        C       D                    �?     ��?             0@        ������������������������       �                     @        E       H                    �?�	j*D�?             *@        F       G                   �a@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        J       O                    b@��S���?             .@       K       L                    @K@      �?              @       ������������������������       �                     @        M       N                   8s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                 ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        S       ^                    �?���@��?            �B@       T       [                   �b@tk~X��?             B@       U       V                    �?��a�n`�?             ?@       ������������������������       �                     9@        W       Z                    �?      �?             @       X       Y                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        \       ]                   `]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        `       �                   @a@.Lj��D�?�             q@       a       �                 pff�?,_ʯ08�?j            �c@       b       i                    �?H%u��?D             Y@        c       d                   �j@     ��?
             0@        ������������������������       �                     @        e       h                   `Y@ףp=
�?             $@        f       g                    �M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        j       o                    �D@(�s���?:             U@        k       n                 ����?�q�q�?             @       l       m                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        p       q                    `@H�!b	�?7            @T@        ������������������������       �                     :@        r       w                    �?,�+�C�?'            �K@        s       v                   �`@z�G�z�?             $@        t       u                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        x       y                    �?`Ӹ����?             �F@        ������������������������       �                     7@        z       �                   @s@�C��2(�?             6@       {       |                    @K@P���Q�?             4@        ������������������������       �                     $@        }       �                    \@ףp=
�?             $@        ~                          �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �_@P����?&            �M@        �       �                   �\@�IєX�?	             1@        �       �                   pp@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     E@        �       �                    @LQI�F�?E            @\@       �       �                 033�?2���?9            �W@       �       �                    �A@:%�[��?*            �Q@        ������������������������       �                     $@        �       �                   �b@N1���?'            �N@       �       �       
             �?��
ц��?"             J@       �       �                   q@�xGZ���?            �A@       �       �                    �?�q�q�?             8@        ������������������������       �                     @        �       �                    �?X�<ݚ�?
             2@       �       �                     E@���Q��?             $@        ������������������������       �                     @        �       �                   @_@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?"pc�
�?	             &@        ������������������������       �                     �?        �       �                   �e@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?�t����?
             1@       �       �                    �?r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        �       �                   �c@���Q��?             @        ������������������������       �                      @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        �       �                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �       	             �?�q�q�?             8@       �       �                    �?�GN�z�?             6@        �       �                    �?�q�q�?             @       �       �                    b@z�G�z�?             @        ������������������������       �                      @        �       �                    c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @e@     ��?             0@        ������������������������       �                     �?        �       �                   �g@�r����?             .@        ������������������������       �                     @        �       �                   �\@"pc�
�?             &@        ������������������������       �                     �?        �       �                   j@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?�X�<ݺ?             2@        ������������������������       �                     "@        �       �                    �G@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��8��,�?g            `c@       �       �       
             �?���tcH�?N            @^@       �       �                    �?�r�MȢ?E            �Z@        �       �                    �M@ףp=
�?             4@        �       �                    �L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �        8            �U@        �       �                    @N@d}h���?	             ,@       ������������������������       �                      @        �       �                   p`@      �?             @        ������������������������       �                      @        �       �                    �N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��.k���?             A@        �       �                    �?      �?             0@        ������������������������       �                     @        �       �                    �Q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �a@r�q��?             2@       �       �                   �`@���!pc�?             &@       �       �                    �?z�G�z�?             $@       �       �                   �^@      �?              @       ������������������������       �                     @        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��C�l�?z?+^���?���S��?���X���?}9�?�F���?�������?�?�䣓�N�?p����?e�kBP��?�	A����?��}A�?�}A_З?�؉�؉�?;�;��?      �?              �?      �?              �?      �?        :�&oe�?�x+�R�?~������?���|?�������?�������?      �?      �?      �?                      �?      �?              �?        ;�;��?;�;��?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?��Hx��?�n���?F]t�E�?t�E]t�?=
ףp=�?
ףp=
�?      �?      �?)\���(�?���Q��?��.���?t�E]t�?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?              �?      �?      �?                      �?      �?        �$I�$I�?�m۶m��?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?��8��8�?�q�q�?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?      �?      �?        ;�;��?vb'vb'�?      �?      �?      �?                      �?              �?�������?�?      �?      �?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        к����?L�Ϻ��?9��8���?r�q��?�c�1Ƹ?�s�9��?              �?      �?      �?      �?      �?      �?                      �?              �?�������?�������?              �?      �?              �?        �������?�������?��J�?����6b�?���Q��?)\���(�?      �?      �?      �?        �������?�������?�������?�������?      �?                      �?              �?��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�����H�?b�2�tk�?              �?��)A��?�}��7��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?l�l��??�>��?              �?F]t�E�?]t�E�?�������?ffffff�?              �?�������?�������?      �?      �?      �?                      �?              �?      �?      �?              �?      �?        'u_[�?�V'u�?�?�?�������?�������?      �?                      �?              �?              �?4��A�/�?f�&_6h�?��=�ĩ�?�a�+�?�'�K=�?+l$Za�?              �?�}�K�`�?�:ڼO�?�;�;�?�؉�؉�?�A�A�?�_�_�?�������?�������?      �?        �q�q�?r�q��?333333�?�������?              �?۶m۶m�?�$I�$I�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?        �������?�������?�������?UUUUUU�?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?UUUUUU�?�������?�袋.��?]t�E�?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?�������?�?      �?        /�袋.�?F]t�E�?              �?�������?�������?              �?      �?              �?        �q�q�?��8��8�?              �?�q�q�?�q�q�?      �?                      �?���/Y��?@��i@�?�C��2(�?����|��?�+J�#�?z����f�?�������?�������?�������?333333�?              �?      �?                      �?              �?۶m۶m�?I�$I�$�?              �?      �?      �?      �?              �?      �?      �?                      �?�������?�?      �?      �?      �?        �q�q�?�q�q�?      �?                      �?UUUUUU�?�������?t�E]t�?F]t�E�?�������?�������?      �?      �?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ �4BhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B@0         f                    �?"�\�&U�?�           ��@               3                    �?01�LՓ�?�            �u@              2                    �R@��8����?�            �j@              	                    \@8�W���?�            `j@                                   �?�z�G��?
             $@                                  �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        
       )                    �? ��A�4�?�             i@              (                   @g@+Rh�r�?z            `g@                                 �c@�g�y��?y            @g@                                  @L@����!p�?>             V@                                 @[@����e��?.            �P@                                   �?�q�q�?             @                                 @q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        +            �O@                                   @N@"pc�
�?             6@                                @33�?      �?             @        ������������������������       �                      @                      
             �?      �?             @        ������������������������       �                      @                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  Pc@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?                '                   e@@uvI��?;            �X@        !       &                   �\@��Y��]�?            �D@        "       %                    �I@z�G�z�?             @        #       $                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        ������������������������       �        %            �L@        ������������������������       �                     �?        *       +                    �?d}h���?             ,@        ������������������������       �                     @        ,       -                 ����?և���X�?             @        ������������������������       �                      @        .       /                    �K@z�G�z�?             @        ������������������������       �                      @        0       1                 ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        4       A                   �a@4;����?W            �`@        5       8                    �?4և����?*             L@        6       7                    �?      �?             0@        ������������������������       �                     @        ������������������������       �                     (@        9       :                   pm@�(\����?             D@       ������������������������       �                     :@        ;       <                    @N@@4և���?
             ,@        ������������������������       �                     @        =       @                    �?      �?              @       >       ?                   �n@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        B       c       	             �?�eP*L��?-            @S@       C       b                   �z@      �?              L@       D       M                     H@r�z-��?            �J@        E       L                   0n@ҳ�wY;�?
             1@       F       K                    �?8�Z$���?             *@       G       J                   �b@�8��8��?             (@        H       I                   @b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        N       W                    �?tk~X��?             B@       O       P                 ����?�����?             5@        ������������������������       �                     �?        Q       R                   �c@P���Q�?             4@       ������������������������       �                     ,@        S       V                    �?r�q��?             @       T       U                 `ff@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        X       a                    �?�q�q�?             .@       Y       `                     P@      �?             $@       Z       [                    �?����X�?             @        ������������������������       �                     �?        \       ]                   �c@r�q��?             @        ������������������������       �                     @        ^       _                   n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        d       e                   p@�q�q�?             5@       ������������������������       �                     ,@        ������������������������       �                     @        g       �                    �?B@!�S3�?�            0x@       h       �                    �?������?�            �r@       i       v                    �?��h#"��?            `j@        j       u                 033�?���"͏�?            �B@       k       r                   �`@8�A�0��?             6@        l       q                    �?z�G�z�?             $@       m       n                   �`@�����H�?             "@       ������������������������       �                     @        o       p                   `]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        s       t                   �u@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �        	             .@        w       z                    �?�w��RR�?h            �e@        x       y                   �W@�t����?             1@        ������������������������       �                      @        ������������������������       �        
             .@        {       �                    �L@�������?]            �c@       |       �                    �?��-#���?=            �Z@        }       �                    �?�n`���?             ?@       ~                           b@�<ݚ�?             ;@        ������������������������       �                     ,@        �       �                   �b@��
ц��?             *@        ������������������������       �                     @        �       �                     E@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �q@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �F@`2U0*��?.            �R@        ������������������������       �                     *@        �       �                    �?Hn�.P��?&             O@       �       �                   �[@�h����?!             L@        �       �                   �a@�IєX�?             1@        �       �                    a@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                    �C@        �       �                   �_@�q�q�?             @       �       �                   �r@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �I@        �       �                    �?���E�?8            �U@        �       �                   �U@��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �        .             R@        �       �                   @E@(����7�?9            @V@        �       �                   �]@      �?             8@        �       �                    �?      �?              @        �       �                    \@z�G�z�?             @        ������������������������       �                      @        �       �                   @Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@      �?             0@       ������������������������       �        	             (@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?؇>���?(            @P@       �       �                    �?�C��2(�?             F@       �       �                   �`@�����H�?             B@        ������������������������       �                     (@        �       �                     N@r�q��?             8@       �       �                   �e@���N8�?             5@       ������������������������       �        
             2@        �       �                    \@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 pff�?և���X�?             5@        �       �                    �?      �?             (@       �       �                    b@      �?              @        �       �                   �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     P@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �t�b�      h�h)h,K ��h.��R�(KK�KK��hi�B  ��j��`�?:�J;�O�?�i#p���?-���?蝺����?�+J�#�?Cs;�G�?��H����?ffffff�?333333�?      �?      �?      �?                      �?              �?��`ph�?�C��x�?͞��X��?*�Ap*�?��{���?�B!��?/�袋.�?]t�E�?�>����?|���?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?        /�袋.�?F]t�E�?      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?      �?                      �?�Cc}h��?9/���?8��18�?������?�������?�������?      �?      �?      �?                      �?      �?              �?              �?                      �?I�$I�$�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�3�τ?�?f�=`�?�m۶m۶?I�$I�$�?      �?      �?      �?                      �?�������?333333�?              �?�$I�$I�?n۶m۶�?              �?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?              �?]t�E�?t�E]t�?      �?      �?�琚`��?����!�?�������?�������?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?              �?9��8���?r�q��?�a�a�?=��<���?      �?        �������?ffffff�?              �?UUUUUU�?�������?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?I��6#�?nF2<��?�1�O
�?�����?��p�C�?�N�с��?*�Y7�"�?v�)�Y7�?/�袋.�?颋.���?�������?�������?�q�q�?�q�q�?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?J��/�?ס�l��?�?<<<<<<�?      �?                      �?b��x�Y�?�fue*�?�琚`��?��sH�?�c�1��?�9�s��?�q�q�?9��8���?              �?�؉�؉�?�;�;�?      �?        �q�q�?9��8���?              �?�������?333333�?              �?      �?                      �?{�G�z�?���Q��?              �?�c�1ƨ?t�9�s�?�$I�$I�?۶m۶m�?�?�?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?Ȥx�L��?m��֡�?�?�������?      �?                      �?              �?<��x��?�9�as�?      �?      �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?      �?      �?                      �?�����? �����?]t�E�?F]t�E�?�q�q�?�q�q�?      �?        �������?UUUUUU�?��y��y�?�a�a�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJڗhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK兔h��B@9         �                    �?&I,|-��?�           ��@                                 �_@h�����?            |@                                   �?��<b���?/            @Q@                                   �?��>4և�?             <@                                  @�d�����?             3@                                  �?�q�q�?	             (@              
                   �\@      �?              @               	                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                   �?�q�q�?             "@                               ����?      �?              @        ������������������������       �                     @                                   �L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                    O@������?            �D@                                  �?@-�_ .�?            �B@                                   �?�<ݚ�?             "@                                  @^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@                                   �?      �?             @       ������������������������       �                      @        ������������������������       �                      @                a                 ����?|��4�5�?�            �w@       !       D                    �?r�q��?�             s@       "       5                    �?�1e�3��?�            �m@       #       $                    �?��e�_�?�            �g@        ������������������������       �        )            �N@        %       0                    @N@     8�?Z             `@       &       '                   �k@P����?R            �]@        ������������������������       �        "             K@        (       )                   @[@      �?0             P@        ������������������������       �                     �?        *       +                    �? ������?/            �O@        ������������������������       �                      @        ,       /                   �k@ �Jj�G�?)            �K@        -       .                   �e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        &             J@        1       2                    �?�z�G��?             $@        ������������������������       �                     @        3       4                     P@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        6       7                    �?��k=.��?            �G@       ������������������������       �                     ?@        8       =                   �q@     ��?
             0@       9       <                    �?      �?              @       :       ;                    \@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        >       ?                    @I@      �?              @        ������������������������       �                     @        @       C                    s@      �?             @       A       B                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        E       X                    �?��(@��?%            �Q@       F       M                     L@�q�q�?            �I@       G       L                   �j@H�V�e��?             A@        H       I                   �f@���|���?             &@        ������������������������       �                     @        J       K                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        N       W                    �?j���� �?
             1@       O       V       	             �?�θ�?             *@       P       S                    �?���!pc�?             &@        Q       R                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                    �O@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Y       Z                 ����?�S����?
             3@        ������������������������       �                     �?        [       \                    @L@�����H�?	             2@       ������������������������       �                     &@        ]       ^                   �`@����X�?             @        ������������������������       �                     �?        _       `                    @N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        b       e                    �?b1<+�C�?*            @R@        c       d                    �?�KM�]�?             3@       ������������������������       �        	             1@        ������������������������       �                      @        f       u                    �?�{��?��?             K@       g       t                    �?     ��?             @@       h       s                 `ff@�E��ӭ�?             2@       i       r                   @b@X�<ݚ�?             "@       j       o                    �?և���X�?             @        k       n       	             �?�q�q�?             @       l       m                   0j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        p       q                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     ,@        v       }                    �?���!pc�?             6@       w       |                    �?r�q��?
             2@       x       {                   �k@���!pc�?             &@        y       z                    @I@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ~                          @l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?T;���?�            �q@        �       �                    �?l��
I��?.            @T@        �       �                   �b@�n_Y�K�?             *@        �       �                    �?����X�?             @       �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@������?&             Q@        �       �                    �?ҳ�wY;�?             A@       �       �                    �?r�q��?             8@       ������������������������       �                     0@        �       �                    �?      �?              @        �       �                   �_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�t����?             A@       �       �                    �?�㙢�c�?             7@        ������������������������       �                     @        �       �                    �?�<ݚ�?             2@       �       �                    _@@�0�!��?
             1@        ������������������������       �                     @        �       �                   �o@      �?             (@       �       �                   `d@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?hL 7Cv�?�            �i@       �       �                    �? ]�� ��?�            �f@        �       �                    �?z�G�z�?             >@       �       �                   pb@8�Z$���?             :@       �       �                    �?���N8�?             5@       �       �                   `c@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �_@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     N@      �?             @        ������������������������       �                     �?        �       �                   Pn@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �R@�.(�i��?k            �b@       �       �                   �U@ "��u�?j            �b@        ������������������������       �                     �?        �       �                   pa@p���?i            �b@       �       �                    �?�?�|�?O            �[@       �       �                    j@�g�y��?C            @W@        �       �                   �h@Du9iH��?            �E@       ������������������������       �                    �A@        �       �                    �?      �?              @       �       �                    �?�q�q�?             @        �       �                    \@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        &             I@        ������������������������       �                     2@        �       �                    �J@�?�'�@�?             C@        �       �                   pk@����X�?	             ,@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             $@        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     N@ �q�q�?             8@       �       �                    c@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?�q�q�?             8@        �       �                    �J@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �X@��
ц��?             *@        �       �                   �_@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?r�q��?             @        �       �                   �e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  �"z?+�?���B`��?�$I�$I�?۶m۶m�?��Moz��?��,d!�?I�$I�$�?۶m۶m�?y�5���?Cy�5��?�������?�������?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?333333�?              �?      �?              �?        ������?�|����?к����?S�n0E�?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?              �?      �?        @��E���?���t	6�?�������?UUUUUU�?�/���?W'u_�?t���G'�?p����?      �?             ��?      �?�V'u�?'u_[�?      �?              �?      �?              �?��}��}�?AA�?      �?        k߰�k�?��)A��?UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?        g���Q��?br1���?      �?              �?      �?      �?      �?�m۶m��?�$I�$I�?              �?      �?              �?              �?      �?              �?      �?      �?      �?      �?              �?      �?                      �?��+��+�?����?UUUUUU�?UUUUUU�?ZZZZZZ�?iiiiii�?]t�E]�?F]t�E�?              �?      �?      �?              �?      �?                      �?�������?ZZZZZZ�?ى�؉��?�؉�؉�?F]t�E�?t�E]t�?      �?      �?      �?                      �?9��8���?�q�q�?      �?                      �?      �?                      �?(������?^Cy�5�?              �?�q�q�?�q�q�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        Ĉ#F��?�;w�ܹ�?�k(���?(�����?      �?                      �?/�����?���^B{�?      �?      �?r�q��?�q�q�?r�q��?�q�q�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?              �?      �?              �?                      �?              �?t�E]t�?F]t�E�?UUUUUU�?�������?t�E]t�?F]t�E�?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?        -)D�{�?�5�n��?h/�����?Lh/����?;�;��?ى�؉��?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?              �?        �?xxxxxx�?�������?�������?UUUUUU�?�������?              �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?        �������?�������?              �?      �?        �?<<<<<<�?d!Y�B�?�7��Mo�?              �?�q�q�?9��8���?�������?ZZZZZZ�?              �?      �?      �?�������?�������?              �?      �?              �?              �?                      �?��߁��?A���@�?�rS�<��?���e�+�?�������?�������?;�;��?;�;��?�a�a�?��y��y�?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?��C�!��?���{��?���Q��?�G�z�?      �?        �3�=l}�?�\"<)H�?к����?*�Y7�"�?�B!��?��{���?w�qGܱ?qG�w��?              �?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?              �?y�5���?������?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?      �?      �?      �?                      �?              �?UUUUUU�?�������?;�;��?�؉�؉�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?F]t�E�?]t�E�?      �?                      �?�;�;�?�؉�؉�?�$I�$I�?�m۶m��?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKÅ�h��B�0         X                    �?�_�6K��?�           ��@                                   �F@�f@���?�            �u@                                  �q@`Ql�R�?4            �W@       ������������������������       �        *            @T@                                  r@8�Z$���?
             *@        ������������������������       �                     �?                                    E@�8��8��?	             (@       ������������������������       �                     $@        	       
       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               E                    �?�j'�]�?�            �o@               2                    �?����3��?G             Z@                                  �?r�q��?2             R@                                  �Z@���B���?             :@                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?�C��2(�?             6@                                   �?�<ݚ�?             "@                                 �g@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                      
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@                                  @\@��+7��?!             G@        ������������������������       �                      @               1                   �e@�����?             C@              "                    �?��R[s�?            �A@                !                 033�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        #       .                    �?r�q��?             >@       $       %       
             �?HP�s��?             9@        ������������������������       �                      @        &       -                    �Q@���}<S�?             7@       '       ,                   @^@���7�?             6@        (       )                   �]@r�q��?             @        ������������������������       �                     @        *       +                   p`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     �?        /       0                   p@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        3       D                 ���@     ��?             @@       4       5                    �?��� ��?             ?@        ������������������������       �                     @        6       =                   @b@؇���X�?             <@       7       <                    @K@P���Q�?             4@        8       9                    �?r�q��?             @        ������������������������       �                     @        :       ;                   ``@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        >       C                   �a@      �?              @       ?       B                    �?���Q��?             @       @       A       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        F       G                    �I@BӀN��?^            �b@        ������������������������       �                     D@        H       Q                    `@���l��?E            �[@        I       P                 @33�?tk~X��?             B@       J       O                   �p@`Jj��?             ?@       K       L                   �a@      �?             0@       ������������������������       �                     &@        M       N                    @L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     @        R       S                 ����?�}��L�?.            �R@       ������������������������       �        $             M@        T       U                    @M@�IєX�?
             1@        ������������������������       �                     (@        V       W                    j@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        Y       �                    �?�ꇗG�?�            x@        Z       �                 ����?`�(c�?_            `b@       [       b                   @E@���>4��?I             \@        \       a                    �?�r����?             >@        ]       `                   �_@����X�?             ,@       ^       _                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        c       t                    �?v�2t5�?8            �T@        d       s                    �?������?             A@       e       j                   �_@     ��?             @@       f       g                 ����?      �?             0@       ������������������������       �        
             ,@        h       i                   Pp@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        k       r                   hq@     ��?
             0@       l       m                    �?�n_Y�K�?             *@        ������������������������       �                     @        n       o                    @K@z�G�z�?             $@        ������������������������       �                     @        p       q                   �l@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        u       �                    �?r�q��?!             H@       v       �                   @b@���y4F�?             C@       w       x                    c@r�q��?             B@        ������������������������       �                     2@        y       z                    \@�q�q�?             2@        ������������������������       �                     @        {       ~                    k@؇���X�?
             ,@        |       }                   Pj@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                   �q@�8��8��?             (@       ������������������������       �                     "@        �       �                    �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?؇���X�?            �A@        �       �                    �?���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                   d@ �q�q�?             8@       ������������������������       �                     6@        �       �                     E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �U@T�W2��?�            �m@        ������������������������       �                     @        �       �                    �? ��Ou��?�            @m@        �       �                    �R@���c���?%             J@       �       �                    �?�t����?$            �I@       �       �                    �?z�G�z�?             >@        ������������������������       �                     �?        �       �                    �?д>��C�?             =@       �       �                   �b@�GN�z�?             6@       �       �                   �`@��s����?             5@        �       �                   0j@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�8��8��?             (@        �       �                    �G@z�G�z�?             @        ������������������������       �                      @        �       �                   �p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                     �?        �       �                   @\@�ȉo(��?f            �f@        �       �                    �M@ףp=
�?             I@       �       �                   �a@д>��C�?             =@       �       �                    @L@�E��ӭ�?
             2@       �       �                    �?     ��?	             0@       �       �                   `[@�8��8��?             (@       ������������������������       �                      @        �       �                    @K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     5@        �       �                   �b@`���i��?H            �`@       �       �                 ����?��d��?A             ^@        �       �                   pb@Pa�	�?            �@@       ������������������������       �                     <@        �       �                   `c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        ,            �U@        �       �                    �?r�q��?             (@       �       �                    q@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  �ԡh6n�?������?4ƚ�?0�甹��?}g���Q�?W�+�ɕ?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?'vb'vb�?��N��N�?UUUUUU�?UUUUUU�?��؉���?ى�؉��?      �?      �?              �?      �?        ]t�E�?F]t�E�?9��8���?�q�q�?۶m۶m�?�$I�$I�?              �?      �?              �?      �?      �?                      �?      �?        Y�B��?zӛ����?              �?^Cy�5�?Q^Cy��?PuPu�?X|�W|��?�������?�������?      �?                      �?UUUUUU�?�������?{�G�z�?q=
ףp�?              �?d!Y�B�?ӛ���7�?F]t�E�?�.�袋�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?      �?        333333�?�������?      �?                      �?      �?              �?      �?�B!��?�{����?              �?�$I�$I�?۶m۶m�?�������?ffffff�?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �7���M�?ـl@6 �?      �?        ��蕱�?5'��Ps�?r�q��?9��8���?���{��?�B!��?      �?      �?      �?        333333�?�������?      �?                      �?      �?                      �?�_,�Œ�?O贁N�?      �?        �?�?      �?        �������?�������?              �?      �?        ���}D�?U����?4և����?������?n۶m۶�?I�$I�$�?�?�������?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?      �?                      �?              �?              �?��+Q��?�ڕ�]��?�?xxxxxx�?      �?      �?      �?      �?              �?      �?      �?              �?      �?              �?      �?ى�؉��?;�;��?      �?        �������?�������?              �?�$I�$I�?�m۶m��?              �?      �?                      �?      �?        �������?UUUUUU�?6��P^C�?(������?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?F]t�E�?]t�E]�?              �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        ��o��o�?MrMr�?      �?        �i�i�?.��-���?�;�;�?;�;��?�?<<<<<<�?�������?�������?      �?        |a���?a���{�?]t�E�?�袋.��?�a�a�?z��y���?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?              �?      �?        h�h��?�~��?�������?�������?|a���?a���{�?r�q��?�q�q�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?                      �?              �?F]t�E�?F]t�E�?�?�������?|���?|���?              �?�������?�������?      �?                      �?              �?UUUUUU�?�������?F]t�E�?]t�E�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�H'jhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�6         N                    �?8}�ý�?�           ��@               +                    @L@��?�            0u@                                  �?�?��,�?�            �m@                                   �?�5��?'             K@                                  @F@�LQ�1	�?!             G@                                   @�t����?             1@              
       	             �?؇���X�?             ,@              	       
             �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                   �K@\-��p�?             =@                                  �?$�q-�?             :@                                  �?`2U0*��?             9@                                   �?ףp=
�?             $@        ������������������������       �                     @                                   �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                ����?      �?              @                                033�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               &                    �?hl �&�?u             g@               %                    @F|/ߨ�?h            @d@       !       $                   @[@@�z�G�?g             d@        "       #                   �Z@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        `            �b@        ������������������������       �                      @        '       (                    @J@�C��2(�?             6@       ������������������������       �                     ,@        )       *                   `e@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ,       C                    �?:�o���?C            @Y@       -       .                 ����?��N`.�?(            �K@        ������������������������       �        
             *@        /       :                    �?և���X�?             E@       0       9                   �r@���Q��?             9@       1       8                   �c@�G��l��?             5@       2       7                   �n@     ��?             0@       3       4                    �?8�Z$���?	             *@       ������������������������       �                     $@        5       6                   @]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ;       @                   @e@@�0�!��?             1@       <       ?                    �?@4և���?             ,@       =       >                   �]@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        A       B       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        D       M                     R@��<b���?             G@       E       H                    �M@؇���X�?             E@        F       G                 @33�?     ��?	             0@       ������������������������       �                     &@        ������������������������       �                     @        I       J                    �? ��WV�?             :@       ������������������������       �                     2@        K       L                 ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        O       �                 ����?p`q�q��?�            �x@        P       �                    �?b��H���?T            �b@       Q       j                    �?X�<ݚ�?=             [@        R       S                    @F@      �?             D@        ������������������������       �                     @        T       Y                    �J@�ʻ����?             A@        U       X                    �F@      �?             (@        V       W                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        Z       c                   �_@���!pc�?             6@       [       \                   �X@8�Z$���?             *@        ������������������������       �                     @        ]       ^                    �?�<ݚ�?             "@        ������������������������       �                     �?        _       b                   �[@      �?              @        `       a                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        d       e                   �`@X�<ݚ�?             "@        ������������������������       �                     @        f       i                    �?r�q��?             @       g       h                     M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        k       |                    �?�������?%             Q@       l       u                    �?~|z����?            �J@        m       n                   �^@�>4և��?             <@        ������������������������       �                     @        o       p                   �c@HP�s��?             9@       ������������������������       �                     1@        q       r                    �?      �?              @        ������������������������       �                     �?        s       t                     J@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        v       w                   @_@z�G�z�?             9@       ������������������������       �                     .@        x       y                    �?      �?             $@        ������������������������       �                     @        z       {                 ����?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        }       ~                    �?�q�q�?             .@        ������������������������       �                     �?               �                     K@X�Cc�?
             ,@        ������������������������       �                     @        �       �                    U@      �?              @        ������������������������       �                     �?        �       �                   �Y@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?             D@        �       �                   `\@      �?             ,@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@        �       �                    _@`Pp�I�?�            �n@        �       �                 033@�<ݚ�?!             K@       �       �                 ��� @�J�4�?              I@       �       �                    �?���y4F�?             C@       �       �                   �U@      �?             @@        ������������������������       �                     �?        �       �                    @Q@��a�n`�?             ?@       �       �                    �?XB���?             =@       �       �                    �?�}�+r��?             3@       �       �                   `_@��S�ۿ?             .@        ������������������������       �                      @        �       �                     H@؇���X�?             @        ������������������������       �                     @        �       �                     M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        �       �                    `@�q�q�?             @       �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �       �                    �?��A� �?v             h@        �       �                    �?r�q��?             E@       �       �                    �?z�G�z�?             >@       �       �                    �?@�0�!��?             1@       �       �                    �?8�Z$���?	             *@       �       �                    �?���Q��?             @       �       �                   0l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                 `ff @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�θ�?
             *@       ������������������������       �                      @        �       �                   ``@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    S@�8��8��?             (@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?P-�T6��?X            �b@       �       �                    c@������?=             \@       �       �                    @J@ �ׁsF�?6             Y@        �       �                    �?(;L]n�?             >@        �       �                   0n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �        %            �Q@        �       �                    �?r�q��?             (@        ������������������������       �                     @        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        �       �                 ����?���Q��?             @        ������������������������       �                     �?        �       �                    a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    Y@$�q-�?            �C@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    @K@      �?             @        ������������������������       �                     �?        �       �                    b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?г�wY;�?             A@        �       �                   �q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     =@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  a[ӿc�?PR Np�?W�m���?R� %�?����?��o��o�?/�����?h/�����?d!Y�B�?Nozӛ��?�������?�������?۶m۶m�?�$I�$I�?9��8���?�q�q�?              �?      �?              �?                      �?�{a���?a����?;�;��?�؉�؉�?{�G�z�?���Q��?�������?�������?              �?�������?�������?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?        ozӛ���?Y�B��?�Hx�5�?�����H�?�������?�������?�������?�������?      �?                      �?      �?                      �?]t�E�?F]t�E�?      �?              �?      �?      �?                      �?�g����?)0��<��?� O	��?��oX���?              �?۶m۶m�?�$I�$I�?333333�?�������?1�0��?��y��y�?      �?      �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �������?ZZZZZZ�?�$I�$I�?n۶m۶�?�������?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?��,d!�?��Moz��?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?O��N���?;�;��?      �?              �?      �?      �?                      �?              �?�3����?
�Z܄�?�|����?�����?�q�q�?r�q��?      �?      �?              �?<<<<<<�?�������?      �?      �?      �?      �?              �?      �?              �?        t�E]t�?F]t�E�?;�;��?;�;��?              �?�q�q�?9��8���?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?r�q��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�?xxxxxx�?�	�[���?��sHM0�?�$I�$I�?�m۶m��?              �?q=
ףp�?{�G�z�?      �?              �?      �?      �?        �m۶m��?�$I�$I�?      �?                      �?�������?�������?              �?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?        UUUUUU�?UUUUUU�?              �?�m۶m��?%I�$I��?              �?      �?      �?              �?�m۶m��?�$I�$I�?              �?      �?        ffffff�?ffffff�?      �?      �?              �?      �?                      �?���2�?.�ݦ���?�q�q�?9��8���?{�G�z�?�z�G��?(������?6��P^C�?      �?      �?      �?        �c�1Ƹ?�s�9��?�{a���?GX�i���?(�����?�5��P�?�?�������?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �LF�W>�?b6�5��?UUUUUU�?�������?�������?�������?�������?ZZZZZZ�?;�;��?;�;��?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?        �؉�؉�?ى�؉��?              �?333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?�`Q�(X�?���t}��?۶m۶m�?I�$I�$�?{�G�z�?�G�z��?�?�������?      �?      �?      �?                      �?              �?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�?�������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�?�������?�������?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��=yhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKх�h��B@4         \                   �`@��}���?�           ��@               %                    �?�L�^�?�            u@                                ����?      �?B             X@                                  ��>����?%             K@        ������������������������       �                      @                      	             �? ��WV�?#             J@                               ����? 	��p�?             =@              	                   �]@`2U0*��?             9@       ������������������������       �        
             0@        
                          0a@�����H�?             "@                                   �?      �?             @        ������������������������       �                      @                                   Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@                                   pb@���N8�?             E@                     	             �?ףp=
�?             >@                                  �? 	��p�?             =@                                 p`@h�����?             <@       ������������������������       �                     7@                                   �?z�G�z�?             @        ������������������������       �                     �?                                  �V@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        !       "                    @N@�q�q�?             (@       ������������������������       �                     @        #       $                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        &       ?                   P`@���K ]�?�             n@        '       8                    �O@ް� ��?E            �Z@       (       7                 ����?���}<S�?=             W@       )       0                   �r@ZՏ�m|�?             �H@       *       /                    �?������?            �D@       +       .                    �?�}�+r��?             C@        ,       -                   �[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     A@        ������������������������       �                     @        1       4                    �?      �?              @        2       3                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       6                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �E@        9       <                    �?�q�q�?             .@       :       ;                    @���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        =       >                   `^@      �?             @       ������������������������       �                      @        ������������������������       �                      @        @       G                    �?��J��i�?U            �`@        A       B                   @l@      �?              @        ������������������������       �                     @        C       D                    �?      �?             @        ������������������������       �                      @        E       F                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        H       W                     Q@ ������?O            �_@       I       V                    �K@`�߻�ɒ?E             [@        J       K                    �?P�Lt�<�?             C@        ������������������������       �                     @        L       U       
             �?      �?             @@       M       N                    �?�g�y��?             ?@        ������������������������       �                      @        O       P                    @K@XB���?             =@       ������������������������       �                     7@        Q       T                   �m@r�q��?             @        R       S                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        +            �Q@        X       Y                    �?�X�<ݺ?
             2@       ������������������������       �                     0@        Z       [                   P`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       �                    �?pw�ت��?�            �x@       ^       a                    I@~�:T��?�            �m@        _       `                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        b       q                   �l@�p����?�            �l@        c       l                    �L@`2U0*��?C             Y@       d       k                   d@�x�E~�?<            @V@        e       j                    �?      �?              @        f       g       
             �?�q�q�?             @        ������������������������       �                     �?        h       i                   Pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        5            @T@        m       p                    @M@"pc�
�?             &@        n       o                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        r       �                   �d@RB)��.�?J             `@       s       ~                    �?������?G            �^@       t       w                    �?X;��?2            @V@        u       v       
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        x       }                   pn@ ��N8�?/             U@        y       z                    n@$�q-�?             *@       ������������������������       �                     &@        {       |                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        '            �Q@               �                   �n@�ʻ����?             A@        �       �                   �^@������?	             .@        ������������������������       �                     @        �       �                   Pb@���|���?             &@        ������������������������       �                     @        �       �                   pe@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   pf@���y4F�?             3@       �       �                   @c@r�q��?             2@        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �H@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?&K�����?`            �c@       �       �                    �?20J�Ws�?X             b@        �       �                   �b@ҳ�wY;�?,             Q@        �       �                   `Y@��� ��?             ?@        ������������������������       �                     �?        �       �                    �?ףp=
�?             >@       �       �                    �?ܷ��?��?             =@        �       �                    a@�q�q�?             @        ������������������������       �                     @        �       �                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 hff�?�nkK�?             7@       ������������������������       �        
             6@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��%��?            �B@       �       �                   �a@`՟�G��?             ?@       �       �                    �?��>4և�?             <@        �       �                   �c@���Q��?	             .@        ������������������������       �                     @        ������������������������       �                     "@        �       �                   Pd@�n_Y�K�?
             *@        �       �                   0j@���Q��?             @        ������������������������       �                      @        �       �                    o@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �V@:���u��?,            @S@        ������������������������       �        	             0@        �       �                    �?�ɞ`s�?#            �N@        �       �                    @K@�G��l��?             5@        �       �                    �F@ףp=
�?             $@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?�C��2(�?             &@        �       �                   �`@z�G�z�?             @        ������������������������       �                      @        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `@R���Q�?             D@        ������������������������       �        
             1@        �       �                    c@�û��|�?             7@       �       �                   �a@������?	             1@       �       �                    �?���Q��?             $@        ������������������������       �                     @        �       �                    b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 033�?r�q��?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B  q��H��?��>���?������?x� O�?      �?      �?�Kh/��?h/�����?              �?O��N���?;�;��?������?�{a���?���Q��?{�G�z�?      �?        �q�q�?�q�q�?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?              �?        ��y��y�?�a�a�?�������?�������?�{a���?������?�$I�$I�?�m۶m��?              �?�������?�������?              �?      �?      �?      �?                      �?      �?              �?        �������?�������?      �?        UUUUUU�?�������?      �?                      �?�N�N�?�,6�,6�?�rp�_��?J�#��?d!Y�B�?ӛ���7�?9/����?�>4և��?������?p>�cp�?(�����?�5��P�?      �?      �?              �?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?�������?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?      �?                      �?      �?      �?              �?      �?        ���@��?�[�՘H�?      �?      �?              �?      �?      �?              �?      �?      �?      �?                      �?AA�?��}��}�?h/�����?B{	�%��?(�����?���k(�?              �?      �?      �?�B!��?��{���?              �?�{a���?GX�i���?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?              �?�q�q�?��8��8�?              �?      �?      �?              �?      �?        Rņ�N�?\u�b��?��7���?@|4!/l�?�������?�������?              �?      �?        T��
��?��e��S�?���Q��?{�G�z�?����G�?p�\��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?        /�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?        S֔5eM�?���)k��?G:l��F�?�On���?�u�{���?�E(B�?333333�?�������?              �?      �?        �y��y��?�a�a�?�؉�؉�?;�;��?      �?              �?      �?              �?      �?              �?        <<<<<<�?�������?wwwwww�?�?      �?        ]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        (������?6��P^C�?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        UUUUUU�?�������?      �?                      �?
�Z܄�?{�ґ=�?�Ő��?z�!���?�������?�������?�{����?�B!��?              �?�������?�������?��=���?a���{�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �Mozӛ�?d!Y�B�?      �?                      �?      �?        }���g�?���L�?�1�c��?�s�9��?۶m۶m�?I�$I�$�?333333�?�������?              �?      �?        ;�;��?ى�؉��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?              �?qV~B���?dj`��?              �?&C��6��?mާ�d�?��y��y�?1�0��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?              �?��,d!�?8��Moz�?�?xxxxxx�?�������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��ChG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B@>         n                 ����?8}�ý�?�           ��@               Y                    �?�LG�4�?�            `v@              P                    �?�șvh�?�            s@              E                    �?�1/z��?�             o@                                  @C@$�� ���?�            �m@                                   �?��X��?             <@              
                    �A@�KM�]�?             3@              	                    �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @                                   �?�<ݚ�?             "@                                  @e@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               :       	             �?(N:!���?�            @j@                                 �a@�i��b��?N            �_@                                  p`@�eP*L��?	             &@                                  �?      �?              @                                  \@      �?             @        ������������������������       �                     �?                                   п�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               #                    �?X�
����?E             ]@                                    �?���|���?             &@                                ����?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        !       "                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        $       1                    @F@����?=            @Z@        %       &                   �h@��+7��?             7@        ������������������������       �                      @        '       .                    �?��s����?             5@       (       -                    @D@�����H�?             2@        )       *                   �f@�<ݚ�?             "@       ������������������������       �                     @        +       ,                   @b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        /       0                   s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        2       3                   �r@��Y��]�?/            �T@       ������������������������       �        )             S@        4       9                   Ps@�q�q�?             @        5       6                   �_@�q�q�?             @        ������������������������       �                     �?        7       8                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ;       <                   `X@P��BNֱ?:            �T@        ������������������������       �                     �?        =       B                   �?��Y��]�?9            �T@       >       A                    �?�(�Tw�?6            �S@       ?       @                   �g@`׀�:M�?3            �R@       ������������������������       �        2            @R@        ������������������������       �                     �?        ������������������������       �                     @        C       D                    �L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        F       O                 ����?�eP*L��?	             &@       G       N                    �?�q�q�?             "@       H       I                   �_@և���X�?             @        ������������������������       �                     �?        J       K                    @A@�q�q�?             @        ������������������������       �                     @        L       M                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        Q       R                   �O@���>4��?             L@        ������������������������       �                     3@        S       X                    �?V������?            �B@        T       U                   �l@�8��8��?             (@       ������������������������       �                     $@        V       W                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        Z       [                    п�c�����?"            �J@        ������������������������       �                     @        \       a                    �?r�qG�?             H@        ]       ^                   �b@�����H�?
             2@       ������������������������       �                     (@        _       `                    �M@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        b       i                    �?d��0u��?             >@        c       h                    h@r�q��?	             (@        d       g                    �?�q�q�?             @       e       f       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        j       k                    p@�X�<ݺ?             2@       ������������������������       �        	             ,@        l       m                    @O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        o       �                   �b@�B!Ae�?�            �w@       p       �                    �?�bW"<�?�            r@       q       �                   {@�]�{���?�            0p@       r       �                   8s@��O���?�            �o@       s       �                    �?�˹�m��?�            �l@        t       y                    �?�q�q�?             H@        u       x                     P@      �?              @       v       w                     M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        z       �                    �?��(\���?             D@        {       �                    �?     ��?
             0@       |       }       
             �?�z�G��?             $@        ������������������������       �                     @        ~                        ����?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        �       �                    �?`Ӹ����?v            �f@       �       �                   @f@г�wY;�?Z             a@        ������������������������       �                    �K@        �       �                    �?H�!b	�?;            @T@        �       �                   �^@؇���X�?
             ,@        ������������������������       �                     @        �       �                   �a@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?0�,���?1            �P@        �       �                   `_@�IєX�?             A@       ������������������������       �                     3@        �       �                    ^@�r����?
             .@        �       �                 ����?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                    �@@        �       �                   �`@�C��2(�?             F@        �       �                   �X@���|���?	             &@        ������������������������       �                     �?        �       �                    �?�z�G��?             $@        ������������������������       �                     �?        �       �                   �]@�q�q�?             "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                   �k@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �@@        �       �                    �?�<ݚ�?             ;@        ������������������������       �                     &@        �       �                    �?      �?	             0@        �       �                    Z@����X�?             @        ������������������������       �                     @        �       �                    ^@�q�q�?             @       �       �                   �v@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @Q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?d��0u��?             >@        �       �                   �a@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?z�G�z�?             4@        �       �                    �?���Q��?             @       �       �                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    `@�r����?
             .@       ������������������������       �                     "@        �       �                    �L@�q�q�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @M@������?6            �U@       �       �                   `T@�q�q�?$             N@        ������������������������       �                     @        �       �                   0a@������?!             K@       �       �                    �?��r._�?            �D@       �       �                    �L@�t����?             A@       �       �                   �f@��S�ۿ?             >@       �       �                   �\@h�����?             <@        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?և���X�?             @       �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �c@��
ц��?             *@        ������������������������       �                      @        �       �                    �?�eP*L��?             &@       �       �                    e@      �?              @       ������������������������       �                     @        �       �                   0m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   c@������?             ;@        ������������������������       �                      @        �       �                    �?z�G�z�?             9@       �       �                   @e@�E��ӭ�?             2@       �       �                   �c@     ��?
             0@       �       �                   y@�z�G��?             $@       �       �                    �?և���X�?             @       �       �                    b@�q�q�?             @       �       �                    �M@      �?             @        ������������������������       �                     �?        �       �                    �N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  a[ӿc�?PR Np�?@aT��A�?=W�l|�?��U���?�+����?��h���?���\V�?l"�k"��?Rv�Qv��?n۶m۶�?%I�$I��?�k(���?(�����?/�袋.�?F]t�E�?      �?                      �?      �?        �q�q�?9��8���?�������?333333�?              �?      �?                      �?|�W|�W�?�A�A�?�V��j��?K�R�T*�?]t�E�?t�E]t�?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        	�=����?���=��?F]t�E�?]t�E]�?333333�?�������?      �?                      �?UUUUUU�?�������?      �?                      �?�؏�؏�?8�8��?zӛ����?Y�B��?              �?z��y���?�a�a�?�q�q�?�q�q�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        8��18�?������?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ��FS���?���ˊ��?              �?8��18�?������?p��o���?�A�A�?��L��?к����?      �?                      �?      �?              �?      �?              �?      �?        ]t�E�?t�E]t�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        n۶m۶�?I�$I�$�?              �?�g�`�|�?o0E>��?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        :�&oe�?�V�9�&�?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?        wwwwww�?DDDDDD�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �q�q�?��8��8�?              �?      �?      �?              �?      �?        �Q�٨��?�+����?��\���?�����?��q/�?�����?�?�������?^Cy�5�?��P^Cy�?�������?UUUUUU�?      �?      �?      �?      �?      �?                      �?      �?        333333�?�������?      �?      �?333333�?ffffff�?              �?333333�?�������?      �?                      �?              �?              �?l�l��??�>��?�?�?              �?�����H�?b�2�tk�?�$I�$I�?۶m۶m�?              �?�$I�$I�?�m۶m��?      �?                      �?g��1��?Ez�rv�?�?�?              �?�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?F]t�E�?]t�E�?F]t�E�?]t�E]�?      �?        333333�?ffffff�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?                      �?�q�q�?9��8���?              �?      �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�q�q�?�q�q�?              �?      �?              �?      �?      �?                      �?wwwwww�?DDDDDD�?ffffff�?333333�?      �?                      �?�������?�������?�������?333333�?      �?      �?              �?      �?              �?        �?�������?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�/�I�?��֡�l�?UUUUUU�?UUUUUU�?              �?B{	�%��?{	�%���?�ڕ�]��?ە�]���?<<<<<<�?�?�������?�?�m۶m��?�$I�$I�?              �?      �?              �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?              �?      �?              �?        �؉�؉�?�;�;�?              �?t�E]t�?]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?{	�%���?B{	�%��?      �?        �������?�������?r�q��?�q�q�?      �?      �?333333�?ffffff�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�y�/hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��B@6         �                    �?8}�ý�?�           ��@              U                   �b@��TE��?           �y@              6                   a@�.*�7�?�            �t@              /                    �?��$���?�            q@              "                   ``@X�aC�U�?�            �m@                                   �?�W�{�5�??            �W@                                   @ >�֕�?            �A@              	                    �?Pa�	�?            �@@        ������������������������       �        
             2@        
                          �q@��S�ۿ?             .@       ������������������������       �                     &@                                    N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                  q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   @L@R���Q�?(             N@                                 �s@�7��?            �C@       ������������������������       �                    �@@                                  �z@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @               !                    �?�q�q�?             5@                                  _@     ��?             0@        ������������������������       �                      @                                   `@      �?              @        ������������������������       �                     @                                   _@z�G�z�?             @       ������������������������       �                     @                                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #       *                    �H@�k~X��?W             b@        $       )                   `c@�X�<ݺ?             2@       %       &                    �F@      �?              @       ������������������������       �                     @        '       (                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        +       ,                   P`@������?L            �_@       ������������������������       �        G             ]@        -       .                   c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        0       5                   �r@�������?             A@       1       2                    �?�n`���?             ?@       ������������������������       �                     0@        3       4                    �?���Q��?             .@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        7       P       	             �?�jTM��?(            �N@       8       A                   �j@r�����?"            �J@        9       >                     L@�q�q�?             2@       :       ;                 033@�����H�?             "@       ������������������������       �                     @        <       =                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ?       @                   b@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        B       C                   0a@(N:!���?            �A@        ������������������������       �                     �?        D       O                    �?l��\��?             A@        E       N                    �?d}h���?             ,@       F       M                    �?      �?             (@       G       H                   �_@�z�G��?             $@        ������������������������       �                     @        I       J                 433�?      �?             @        ������������������������       �                     �?        K       L                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     4@        Q       R                    �?      �?              @        ������������������������       �                     �?        S       T                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        V       s                    �?V�K/��?4            �S@       W       ^                    �?x�K��?!            �I@        X       Y                    �?���7�?             6@       ������������������������       �                     .@        Z       [                   0m@؇���X�?             @       ������������������������       �                     @        \       ]                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       d                    �?J�8���?             =@        `       c                   e@z�G�z�?             @        a       b                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        e       j                    @E@      �?             8@        f       i                    @      �?              @       g       h                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        k       r                    �?      �?
             0@       l       q                    �?��S�ۿ?	             .@        m       n                 ����?z�G�z�?             @        ������������������������       �                      @        o       p                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        t       �                    �?d}h���?             <@       u       �                   �r@      �?             0@       v       y                    �?�θ�?
             *@        w       x                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        z       {                     I@      �?              @        ������������������������       �                     @        |                          �c@�q�q�?             @       }       ~                    @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �       	             �?�l8ɠ��?�            t@       �       �                   �`@3�E�?�             j@        �       �                    �?~h����?"             L@       �       �                   �U@p9W��S�?             C@        ������������������������       �                      @        �       �                   `c@      �?             B@       �       �                   �?\-��p�?             =@       ������������������������       �                     2@        �       �                   �U@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                    X@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�����H�?             2@       ������������������������       �                     *@        �       �                 033�?���Q��?             @        ������������������������       �                      @        �       �                    @N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@���y4F�?a             c@       �       �                    �?��0{9�?]            �a@       �       �                 ���ٿ��Ns��?P            �^@        ������������������������       �                     @        �       �       
             �?0y����?O            �]@       �       �                    �?�GN�z�?+            �P@       �       �                    �?d}h���?#             L@        �       �                 033�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @E@z�G�z�?             I@        ������������������������       �                     �?        �       �                    �M@Jm_!'1�?            �H@       �       �                   �c@�ݜ�?            �C@        ������������������������       �        	             (@        �       �                    �D@�+$�jP�?             ;@        �       �                   �\@      �?             @        ������������������������       �                     �?        �       �                    @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �_@�LQ�1	�?             7@        �       �                   Pq@���!pc�?             &@       �       �                   pe@z�G�z�?             $@        �       �                   pd@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   @d@���Q��?             $@       �       �                   �b@և���X�?             @       �       �                   �n@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `m@�z�G��?             $@        ������������������������       �                     @        �       �                 ����?���Q��?             @       �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    c@�O4R���?$            �J@        �       �                   �b@ �q�q�?             8@       ������������������������       �                     7@        ������������������������       �                     �?        ������������������������       �                     =@        �       �                   �Y@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     &@        �       �                    �?���͡?G            @\@        ������������������������       �                     :@        �       �                   �a@�d���?8            �U@        �       �                   �_@`Jj��?             ?@        �       �                   (p@      �?              @        ������������������������       �                     @        �       �                    �K@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     7@        ������������������������       �        %             L@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  a[ӿc�?PR Np�?-m�C��?���/D�?ՃF��[�?�/7Āt�?J�J��?��k��k�?Tn�wp٫?���hB�?Fڱa��?�ĩ�sK�?�A�A�?��+��+�?|���?|���?              �?�?�������?              �?      �?      �?              �?      �?              �?      �?      �?                      �?333333�?333333�?�A�A�?��[��[�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?        �������?�������?      �?              �?      �?      �?                      �?              �?�q�q�?�8��8��?�q�q�?��8��8�?      �?      �?              �?      �?      �?              �?      �?                      �?AA�?�������?              �?�������?�������?              �?      �?        �������?�������?�c�1��?�9�s��?              �?�������?333333�?      �?                      �?      �?        .�u�y�?�y��!�?�V�9�&�?Dj��V��?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?r�q��?�q�q�?      �?                      �?�A�A�?|�W|�W�?      �?        �������?------�?۶m۶m�?I�$I�$�?      �?      �?333333�?ffffff�?              �?      �?      �?      �?        �������?333333�?      �?                      �?              �?              �?              �?      �?      �?              �?�m۶m��?�$I�$I�?      �?                      �?�Z܄��?�ґ=�?ssssss�?�?�.�袋�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?|a���?�rO#,��?�������?�������?      �?      �?              �?      �?              �?              �?      �?      �?      �?�������?UUUUUU�?      �?                      �?              �?      �?      �?�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?۶m۶m�?I�$I�$�?      �?      �?�؉�؉�?ى�؉��?�������?�������?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?���C��?����R�?�N��N��?vb'vb'�?%I�$I��?�m۶m��?�k(����?l(�����?              �?      �?      �?a����?�{a���?      �?        ]t�E]�?F]t�E�?              �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?�q�q�?�q�q�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?6��P^C�?(������?m�w6�;�?L� &W�?7�S\2�?&C��6��?              �?�������?�5�5�?�袋.��?]t�E�?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?����X�?������?\��[���?�i�i�?      �?        /�����?B{	�%��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?��Moz��?Y�B��?F]t�E�?t�E]t�?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        333333�?�������?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?        ffffff�?333333�?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?:�&oe�?�x+�R�?�������?UUUUUU�?      �?                      �?      �?        �k(���?(�����?              �?      �?                      �?$��Co�?x�!���?      �?        �:���C�?Ȥx�L��?���{��?�B!��?      �?      �?      �?        333333�?�������?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�-4FhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK˅�h��B�2         |                    �?6������?�           ��@                               ����?�����?            y@                                   �?��`qM|�?4            �T@                      	             �?ȵHPS!�?             :@                                  �?R���Q�?             4@                                  �?z�G�z�?             .@                                 @b@�z�G��?             $@       ������������������������       �                     @        	       
                    �F@      �?             @        ������������������������       �                      @                                  pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                   �?0�)AU��?#            �L@       ������������������������       �                     H@                                    I@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @               {                    �R@T��ٟK�?�            �s@              F                    �?��t���?�            �s@               !                 pff�?Fx$(�??             Y@                                  @l@؇���X�?             ,@        ������������������������       �                     @                                    �?      �?              @                               ����?�q�q�?             @                      	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        "       E                   @f@�^�����?4            �U@       #       *                    �?rEC��a�?1            �S@        $       %                   `X@�����?             3@        ������������������������       �                      @        &       )                    `P@������?
             1@       '       (                    �?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        +       @                    �?ףp=
�?&             N@       ,       1                    �?�+$�jP�?             ;@        -       0                    �?�q�q�?             @       .       /                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        2       ?                   �n@؇���X�?             5@       3       <                    �?      �?             (@       4       5                   0b@z�G�z�?	             $@        ������������������������       �                     @        6       7                    �K@�q�q�?             @        ������������������������       �                     @        8       9       
             �?�q�q�?             @        ������������������������       �                     �?        :       ;                   d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        =       >                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        A       B                    �?Pa�	�?            �@@       ������������������������       �                     >@        C       D                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        G       `                   �`@�8��8��?�             k@       H       _                    �? ��WV�?g            �c@       I       ^                    �? ѯ��?H            �Z@       J       S                 ����?�*v��?@            @X@        K       R                   �`@�q�q�?             8@       L       M                   �o@X�Cc�?
             ,@        ������������������������       �                     @        N       O                    `@����X�?             @        ������������������������       �                     @        P       Q       
             �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        T       U                 ���@ �й���?/            @R@       ������������������������       �        &             L@        V       ]                   �\@�IєX�?	             1@       W       \                    @�����H�?             "@       X       Y                   �Z@      �?              @        ������������������������       �                     @        Z       [                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                    �H@        a       l                   �j@z�G�z�?'             N@        b       c                    �?�G�z��?             4@        ������������������������       �                     @        d       e                    �?������?             .@        ������������������������       �                     @        f       g                    �?X�<ݚ�?             "@        ������������������������       �                     @        h       k                    �H@r�q��?             @        i       j                   �g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        m       t       
             �?��(\���?             D@       n       o                    @M@�g�y��?             ?@       ������������������������       �                     5@        p       s                     N@ףp=
�?             $@        q       r                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        u       x                    �?�<ݚ�?             "@        v       w                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        y       z                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        }       �                    �?b:�&���?�            �t@       ~       �                    �?L��B�?�            �q@               �                   @c@��<b�ƥ?3             W@       ������������������������       �        .            �U@        �       �                    �?�q�q�?             @       �       �                   �r@z�G�z�?             @        ������������������������       �                     @        �       �                    @O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �O@�m	{�?r            �g@        �       �                   �[@���Q��?             4@        ������������������������       �                     @        �       �                   @^@և���X�?	             ,@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	             �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�� ND��?f            `e@       �       �                    �?���(-�?V            @b@       �       �                   �t@�8���?G             ]@       �       �                    �?�nkK�?F            �\@       �       �                   �? pƵHP�?A             Z@       �       �                    �?�q�q�?:             X@       �       �       	             �?��'�`�?3            �T@        �       �                 ����?�?�|�?            �B@       �       �                   �c@��?^�k�?            �A@        �       �                   �]@      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     3@        ������������������������       �                      @        ������������������������       �                     G@        ������������������������       �                     *@        �       �                   p`@      �?              @        �       �                   �^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pp@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        �       �                   0b@���Q��?             9@        ������������������������       �                      @        �       �                    �?j���� �?             1@       �       �                    �H@�z�G��?             $@        ������������������������       �                     @        �       �                    e@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �P@`�(c�?            �H@       �       �       
             �?�X����?             F@       �       �                    �?�^�����?            �E@       �       �                    �I@�q�q�?             >@        �       �                   Pj@�q�q�?             (@        �       �                 033�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �e@�����H�?             2@       �       �                   �q@�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     M@�θ�?             *@        ������������������������       �                      @        �       �                    S@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��X�5�?��S�$e�?\�՘H�?���-��?��k���?�@	o4u�?�؉�؉�?��N��N�?333333�?333333�?�������?�������?333333�?ffffff�?              �?      �?      �?      �?              �?      �?      �?                      �?              �?              �?              �?p�}��?��Gp�?              �?�q�q�?�q�q�?      �?                      �?�k���?e�}��?^-n����?�td�@T�?R���Q�?ףp=
��?۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ֔5eMY�?�5eMYS�?�=Q���?�0���M�?Q^Cy��?^Cy�5�?              �?xxxxxx�?�?333333�?�������?      �?                      �?      �?        �������?�������?B{	�%��?/�����?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?              �?|���?|���?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?;�;��?O��N���?�@�Ե�?n���4�? tT����?���AG�?�������?UUUUUU�?�m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?                      �?����?����Ǐ�?              �?�?�?�q�q�?�q�q�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?              �?�������?�������?�������?�������?      �?        �?wwwwww�?              �?�q�q�?r�q��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?333333�?�������?�B!��?��{���?              �?�������?�������?�������?�������?              �?      �?                      �?�q�q�?9��8���?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?        �b��7�?o4u~�!�?��/���?�s�vG#�?��7��M�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?                      �?�h�O�?�]Ɣ���?�������?333333�?              �?�$I�$I�?۶m۶m�?۶m۶m�?�$I�$I�?      �?                      �?�$I�$I�?�m۶m��?              �?      �?        �_@�?@���?��իW��?�P�B�
�?j��FX�?a���{�?�Mozӛ�?d!Y�B�?'vb'vb�?;�;��?�������?UUUUUU�?1P�M��?��k���?*�Y7�"�?к����?_�_��?�A�A�?      �?      �?              �?      �?              �?              �?              �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        F]t�E�?t�E]t�?      �?                      �?              �?      �?        333333�?�������?      �?        ZZZZZZ�?�������?ffffff�?333333�?      �?        �������?333333�?      �?                      �?              �?4և����?������?]t�E]�?�E]t��?֔5eMY�?�5eMYS�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?                      �?�q�q�?�q�q�?�?�?              �?      �?              �?        �؉�؉�?ى�؉��?              �?333333�?�������?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJr��<hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKㅔh��B�8         �                    �?�#i����?�           ��@              Q                    �?L�o���?           P{@              >                 ����?�yk�~��?�            s@              =                   h@�<_���?�             q@                                  U@$�q-�?�            q@                                  �R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	                          @E@0M����?�            �p@        
                           �?�E��ӭ�?             2@                                  �?�r����?
             .@                                  �?r�q��?	             (@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?ףp=
�?             $@        ������������������������       �                     @                                    F@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               0                    @L@���T��?�            �o@              +                 ����?�k��$�?x            `h@                                   �?hl �&�?r             g@                                 @[@�k.s�׌?[            �a@                                   �?؇���X�?             @       ������������������������       �                     @                      	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        V            �`@        !       *                    �?X�EQ]N�?            �E@       "       '                    �?r�q��?             >@       #       &                 ����?$�q-�?             :@       $       %                   �b@���}<S�?             7@       ������������������������       �                     5@        ������������������������       �                      @        ������������������������       �                     @        (       )                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        ,       -                    �?"pc�
�?             &@       ������������������������       �                     @        .       /                 ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        1       <                    �?�y��*�?!             M@       2       3                   �n@؇���X�?            �H@       ������������������������       �                     >@        4       ;                   pe@p�ݯ��?             3@       5       :                    �?��S���?             .@       6       9                   �q@�q�q�?             (@        7       8                     O@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ?       F                    �M@���@M^�?             ?@       @       A                    `@j���� �?             1@        ������������������������       �                     @        B       C                 ���@�C��2(�?             &@       ������������������������       �                     @        D       E                 ���
@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        G       P       
             �?؇���X�?	             ,@       H       I                   �^@�<ݚ�?             "@        ������������������������       �                     @        J       M                    �?���Q��?             @       K       L                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        N       O                    @O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        R       �       	             �?�F.< �?V            �`@       S       n                    �? ��(��?K            @\@       T       _                    �?�̨�`<�?9            @U@        U       V                    �D@�q�q�?
             (@        ������������������������       �                     @        W       X                     H@X�<ݚ�?	             "@        ������������������������       �                     @        Y       ^                    �?�q�q�?             @       Z       ]       
             �?z�G�z�?             @       [       \                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        `       m                   �r@F��}��?/            @R@       a       l                    �? �q�q�?.             R@       b       i                    @M@t��ճC�?             F@       c       d                   0a@��Y��]�?            �D@       ������������������������       �                     ;@        e       f                 ����?@4և���?             ,@        ������������������������       �                     "@        g       h                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        j       k                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     <@        ������������������������       �                     �?        o       t                    �?��>4և�?             <@        p       s                    �O@�<ݚ�?             "@        q       r                    @L@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        u       �                   @d@���y4F�?             3@       v       {                    �?�t����?
             1@       w       z                    W@$�q-�?             *@        x       y                    �P@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        |       }                   �c@      �?             @        ������������������������       �                      @        ~                        ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �^@D�n�3�?             3@        �       �                    �I@�����H�?             "@        �       �                     D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @K@F�����?�            �r@        �       �                   �b@ڍ`�ڴ�?B            �\@       �       �                    �?�"�q��?7            �W@        �       �                    �?�q�q�?             (@       �       �                 033�?���!pc�?             &@       �       �                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?��Lɿ��?/            �T@        �       �                    �?�n_Y�K�?             *@        ������������������������       �                      @        �       �                    �I@�eP*L��?             &@       �       �                   �s@      �?              @       �       �                    @D@؇���X�?             @        ������������������������       �                      @        �       �                 ����?z�G�z�?             @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pa@ >�֕�?'            �Q@       �       �                    @J@��v$���?"            �N@       ������������������������       �                    �H@        �       �                    �J@�8��8��?             (@        �       �                    �?r�q��?             @       �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             "@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?             4@        ������������������������       �                     @        �       �                    �?     ��?	             0@        �       �                    �?�z�G��?             $@       �       �                   `e@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �e@�q�q�?             @       �       �                   0k@�q�q�?             @        ������������������������       �                     �?        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   0h@���'\�?s            �f@        �       �                    �?���J��?"            �I@       ������������������������       �                    �C@        �       �                   @b@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �[@A5Xo�?Q            ``@        �       �                   �a@��
ц��?             *@       �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        �       �                   �p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? ,��-�?J            �]@        �       �                   �_@z�G�z�?             4@       ������������������������       �        	             &@        �       �                    �?X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@@9G��?<            �X@       �       �                    �?l�b�G��?"            �L@       �       �                    �?Du9iH��?            �E@        �       �                   �r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?P���Q�?             D@        �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     A@        �       �                    @N@@4և���?	             ,@        ������������������������       �                     @        �       �                     O@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        �t�b�      h�h)h,K ��h.��R�(KK�KK��hi�B0  �5�;���?%e��?u�	���?�����?�4��ǲ�?|,���4�?p�h�?n�?ܺ���?�؉�؉�?;�;��?      �?      �?      �?                      �?��z�l��?��)��?�q�q�?r�q��?�������?�?�������?UUUUUU�?      �?      �?              �?      �?        �������?�������?      �?        �������?UUUUUU�?              �?      �?              �?                      �?�R��N�?qК3[�?�����?PP�?ozӛ���?Y�B��?"����?t�n��}?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        w�qG�?qG�wĽ?�������?UUUUUU�?�؉�؉�?;�;��?ӛ���7�?d!Y�B�?      �?                      �?      �?              �?      �?              �?      �?              �?        /�袋.�?F]t�E�?      �?              �?      �?              �?      �?        �4�rO#�?GX�i��?۶m۶m�?�$I�$I�?      �?        ^Cy�5�?Cy�5��?�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?              �?                      �?      �?              �?                      �?�c�1��?�s�9��?�������?ZZZZZZ�?              �?]t�E�?F]t�E�?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?�q�q�?9��8���?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?                      �?>����?|��|�?Vzja���?ja��V�?�?�������?�������?�������?              �?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ����?��Ǐ?�?UUUUUU�?�������?t�E]t�?�E]t��?������?8��18�?              �?�$I�$I�?n۶m۶�?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        I�$I�$�?۶m۶m�?9��8���?�q�q�?      �?      �?      �?                      �?      �?        (������?6��P^C�?�?<<<<<<�?;�;��?�؉�؉�?�������?�������?              �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?              �?        l(�����?(������?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        ^[�'�A�?)iv���?�����?r�.�|�?|n�S���?a�+F�?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?�q�q�?�q�q�?              �?      �?                      �?              �?rY1P»?�������?ى�؉��?;�;��?              �?]t�E�?t�E]t�?      �?      �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?      �?                      �?              �?      �?              �?        �A�A�?��+��+�?;ڼOqɐ?.�u�y�?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?      �?              �?      �?ffffff�?333333�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        �Q�Q�?��\��\�?�?______�?              �?UUUUUU�?UUUUUU�?              �?      �?        #����[�?��℔�?�؉�؉�?�;�;�?�q�q�?9��8���?              �?      �?      �?      �?                      �?      �?        'u_[�?[4���?�������?�������?              �?�q�q�?r�q��?              �?      �?        9/���?������?p�}��?�Gp��?w�qGܱ?qG�w��?UUUUUU�?UUUUUU�?              �?      �?        �������?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�D�thG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         j                    �?znt��s�?�           ��@               -                    �K@R�|[��?�            `w@              "                 033�? ���x�?�            @l@                                  �?�IJ��?�            @j@                               ���ٿ��?}�?o             g@        ������������������������       �                     �?                                   �?��3EaǼ?n             g@              	                    �?PÅ�R1�?k            �f@       ������������������������       �        O            �`@        
                           @D@Jm_!'1�?            �H@                                   �?      �?             $@        ������������������������       �                     �?                                  �a@X�<ݚ�?             "@                                 �Z@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?��-�=��?            �C@                                 �_@�8��8��?             B@                                ����?      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     8@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   ^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?               !                   @\@ �o_��?             9@                                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        #       $                    �?     ��?             0@        ������������������������       �                     @        %       &                   `T@X�<ݚ�?             "@        ������������������������       �                     @        '       ,                    p@r�q��?             @       (       +                    �I@�q�q�?             @       )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        .       Y                    �?r�J���?U            �b@       /       X                    �R@8^s]e�?0            �U@       0       M                 `ff�?�t����?/            @U@       1       F       	             �?�'�`d�?#            �P@       2       E                   0d@�*/�8V�?            �G@       3       D                   �u@^������?            �A@       4       A                 ����?�f7�z�?             =@       5       :       
             �?�G�z��?             4@       6       9                   �`@�n_Y�K�?             *@       7       8                   �X@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ;       @                   �b@և���X�?             @       <       =                   @^@z�G�z�?             @        ������������������������       �                      @        >       ?                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        B       C                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        G       H                   �a@�KM�]�?             3@        ������������������������       �                     "@        I       J                    @L@z�G�z�?             $@        ������������������������       �                     @        K       L                    �L@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        N       W                   @o@D�n�3�?             3@       O       R                 ����?��S���?
             .@        P       Q                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        S       T                    �?�<ݚ�?             "@        ������������������������       �                     @        U       V                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Z       e                    �?�jTM��?%            �N@       [       `                 033�?���@M^�?             ?@       \       ]                    �L@�\��N��?             3@        ������������������������       �                     @        ^       _                    �?      �?	             (@        ������������������������       �                     @        ������������������������       �                     "@        a       d                    �M@r�q��?             (@        b       c                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        f       i                    @ףp=
�?             >@        g       h                    �R@@�0�!��?             1@       ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �        	             *@        k       �                   �b@�r����?�            �v@       l       �                    �?l'��`�?�            �s@        m       x                    `@tk~X��?1             R@       n       w                    �?�8��8��?             B@        o       t                    �P@�z�G��?	             $@       p       s                    �L@؇���X�?             @        q       r                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        u       v                    k@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        y       �                   �d@<ݚ)�?             B@       z       �                    �?����X�?            �A@       {       �                 hff�?���Q��?             9@        |                           �F@�θ�?             *@        }       ~                     C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     J@�q�q�?             (@        �       �                   �`@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �]@@:��JU�?�            @n@        �       �                   `[@���1��?@            �Z@       ������������������������       �        %            @P@        �       �                    �?�Ń��̧?             E@       �       �                    �L@      �?             @@       �       �                    �?      �?
             0@       �       �                    �?$�q-�?             *@        �       �                    @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     $@        �       �                    �?���?S            �`@        �       �                    �?���y4F�?             3@       �       �                    �?�r����?	             .@       �       �                   �_@$�q-�?             *@        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �s@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 `ff�?XB���?H             ]@       �       �                   `_@�L#���?*            �P@        ������������������������       �                     <@        �       �                 033�?��-�=��?            �C@       �       �                   �l@г�wY;�?             A@       ������������������������       �                     6@        �       �                    �?�8��8��?             (@       �       �                    �?ףp=
�?             $@        �       �                   �n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    Y@���Q��?             @        ������������������������       �                     �?        �       �                   @_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �H@        �       �                    �?(옄��?!             G@        �       �                    �?     ��?             0@       �       �                    �L@$�q-�?	             *@       ������������������������       �                     $@        �       �                   @^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   ``@�q�q�?             @        ������������������������       �                     �?        �       �                   Pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���Q��?             >@       �       �                    �D@�G��l��?             5@        ������������������������       �                     "@        �       �       	             �?�8��8��?             (@       �       �                 ����?�C��2(�?             &@        �       �                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �       
             �?�����H�?             "@       �       �                     K@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  ����?��}t��?0G��/�?�q��+��?	�����?��	���?�����?�r)�r)�?��ׄ���?�	A����?              �?!Y�B�?�Mozӛ�?�!H��h�?��}kdu�?      �?        ����X�?������?      �?      �?      �?        �q�q�?r�q��?�������?�������?              �?      �?                      �?}˷|˷�?�A�A�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        
ףp=
�?�Q����?�q�q�?9��8���?      �?                      �?      �?              �?      �?              �?r�q��?�q�q�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        v�)�Y7�?��L��?|a���?	�=����?�������?�������?6�d�M6�?'�l��&�?�٨�l��?AL� &W�?uPuP�?_�_��?O#,�4��?a���{�?�������?�������?ى�؉��?;�;��?�m۶m��?�$I�$I�?              �?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?�q�q�?      �?                      �?      �?              �?        �k(���?(�����?      �?        �������?�������?      �?        333333�?�������?              �?      �?        (������?l(�����?�?�������?UUUUUU�?�������?      �?                      �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?.�u�y�?�y��!�?�c�1��?�s�9��?y�5���?�5��P�?      �?              �?      �?      �?                      �?UUUUUU�?�������?�������?333333�?      �?                      �?              �?�������?�������?�������?ZZZZZZ�?              �?      �?                      �?�?�������?��O[h��?C����?9��8���?r�q��?UUUUUU�?UUUUUU�?333333�?ffffff�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�8��8��?��8��8�?�$I�$I�?�m۶m��?�������?333333�?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?�������?�������?�$I�$I�?�m۶m��?      �?                      �?      �?                      �?      �?        "pc�
�?��i�V��?�+J�#�?�S�rp��?              �?�a�a�?��<��<�?      �?      �?      �?      �?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?              �?              �?              �?t��:W�?��oS��?(������?6��P^C�?�?�������?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?      �?      �?                      �?�{a���?GX�i���?g��1��?��@���?              �?�A�A�?}˷|˷�?�?�?              �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?333333�?�������?              �?      �?      �?      �?                      �?              �?���,d�?ӛ���7�?      �?      �?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?333333�?1�0��?��y��y�?              �?UUUUUU�?UUUUUU�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?        �q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�o7hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�7         �                    �?0����?�           ��@              %                    �?.P�'z�?           `{@                                   �?\��_��?-            �Q@                                  �?b�2�tk�?             B@        ������������������������       �                     @                                   \@�q�q�?            �@@        ������������������������       �                     @                                  �b@������?             >@       	                           �?8�Z$���?             :@       
                           �?�nkK�?             7@       ������������������������       �                     0@                                   �?؇���X�?             @        ������������������������       �                     @                                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               "                    �?">�֕�?            �A@                                  �?���B���?             :@        ������������������������       �                     @                                   �J@      �?             4@                                   �G@      �?              @        ������������������������       �                     @                                ����?z�G�z�?             @        ������������������������       �                     @                                  Pn@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               !                    �?�8��8��?
             (@                                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        #       $                    �I@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        &       i       
             �?0<o�Ɲ�?�            �v@       '       `       	             �?p���p�?�            Ps@       (       /                    �?�x�+���?�            @r@        )       *                 ����?z�G�z�?             9@        ������������������������       �                     (@        +       .                   �l@�n_Y�K�?             *@        ,       -                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        0       K                 ����?�{��?�            �p@        1       4                   �Q@\#r��?G            �^@        2       3                   �l@      �?             @        ������������������������       �                     @        ������������������������       �                     @        5       6                 ����?,Z0R�?E             ]@        ������������������������       �        !            �J@        7       8                 833�?؇���X�?$            �O@        ������������������������       �                     �?        9       B                 `ff�?��� ��?#             O@        :       A                    �?l��\��?             A@       ;       <                    �?R���Q�?             4@        ������������������������       �                     @        =       @                   `c@     ��?
             0@       >       ?                   �i@�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        C       J                    �?�>4և��?             <@        D       E                   �Y@�n_Y�K�?             *@       ������������������������       �                     @        F       I                   �]@r�q��?             @       G       H                   (q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        L       _                    �?XB���?[             b@       M       T                   `P@��	,UP�?>             W@        N       S                   P`@�<ݚ�?             "@       O       P                    �?      �?              @       ������������������������       �                     @        Q       R                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        U       X                 ����?P��BNֱ?8            �T@        V       W                   �p@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        Y       \                    �?�?�|�?3            �R@       Z       [                   �b@ �Jj�G�?&            �K@       ������������������������       �        %             K@        ������������������������       �                     �?        ]       ^                   �Z@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                    �J@        a       h                    �?��.k���?             1@       b       c                   @`@���Q��?
             .@        ������������������������       �                     @        d       e                    @C@���Q��?             $@        ������������������������       �                     @        f       g                    @L@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        j       w                   �`@T����1�?$             M@        k       r                   �c@�r����?             >@       l       q                   P`@ �q�q�?             8@        m       n                    �?�����H�?             "@       ������������������������       �                     @        o       p                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        s       v                   `Z@      �?             @        t       u                   @W@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        x       �                    �?���>4��?             <@       y       �                    b@\X��t�?             7@       z       �                    �?�����?             3@       {       �                 `ff@�	j*D�?	             *@       |       �                    @N@      �?             (@       }       ~                    �?ףp=
�?             $@       ������������������������       �                      @               �                   m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �k@�q�q�?             @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @E@|��+�?�            �r@        �       �       	             �?��+7��?             7@       �       �                   �?R���Q�?             4@        �       �                   �_@�q�q�?             @        ������������������������       �                     @        �       �                    @O@�q�q�?             @       �       �                   Pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@4և���?
             ,@       �       �                   @`@      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@���f�K�?�            q@       �       �                   �g@ ��� �?�            �j@       �       �                    @D@ 5x ��?�            �j@        �       �                    �?��(\���?             D@       ������������������������       �                    �A@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����? _�@�Y�?j            �e@       �       �                 ����?��f�{��?h            �e@       �       �                    @F@�=
ףp�?_             d@        �       �                   xq@������?             B@       ������������������������       �                     =@        �       �                   (r@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        G             _@        �       �                   �j@�8��8��?	             (@        �       �                   pi@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?8^s]e�?(             M@       �       �                   `]@@�0�!��?             A@        ������������������������       �                      @        �       �                 033@      �?             @@       �       �                   �c@��a�n`�?             ?@        ������������������������       �                     �?        �       �                    �?��S�ۿ?             >@       �       �                   �? ��WV�?             :@       ������������������������       �        
             *@        �       �                   p@$�q-�?             *@       ������������������������       �                     $@        �       �                 pff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@      �?             @        ������������������������       �                      @        �       �                    h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �R@      �?             8@       �       �                   �`@���Q��?             4@        �       �                   �p@�q�q�?             "@       �       �                 ����?      �?             @        ������������������������       �                      @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?"pc�
�?	             &@       �       �                   @l@      �?              @        ������������������������       �                     �?        �       �       
             �?؇���X�?             @       �       �                   �b@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ���^L�?���Y�?j�����?%���V�?�K=��?$Zas �?�8��8��?9��8���?              �?UUUUUU�?UUUUUU�?              �?wwwwww�?�?;�;��?;�;��?�Mozӛ�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?              �?�A�A�?_�_��?ى�؉��?��؉���?              �?      �?      �?      �?      �?              �?�������?�������?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?%e��?���>��?C��ڸ?�E|���?�4iҤI�?mٲe˖�?�������?�������?              �?ى�؉��?;�;��?�m۶m��?�$I�$I�?      �?                      �?              �?�2A�L�?ߥ�wi��?XG��).�?��:��?      �?      �?              �?      �?        	�=��ܳ?�FX�i��?              �?�$I�$I�?۶m۶m�?      �?        �B!��?�{����?�������?------�?333333�?333333�?              �?      �?      �?�?�������?              �?      �?              �?                      �?�m۶m��?�$I�$I�?ى�؉��?;�;��?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�{a���?GX�i���?��Mozӫ?d!Y�B�?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ���ˊ��?��FS���?�q�q�?�q�q�?              �?      �?        к����?*�Y7�"�?��)A��?k߰�k�?              �?      �?        (�����?�5��P�?      �?                      �?              �?�?�������?�������?333333�?              �?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?        �rO#,��?�FX�i��?�?�������?UUUUUU�?�������?�q�q�?�q�q�?              �?      �?      �?      �?                      �?              �?      �?      �?      �?      �?              �?      �?                      �?I�$I�$�?n۶m۶�?��Moz��?!Y�B�?^Cy�5�?Q^Cy��?;�;��?vb'vb'�?      �?      �?�������?�������?              �?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        Z7�"�u�?�"�u�)�?Y�B��?zӛ����?333333�?333333�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �$I�$I�?n۶m۶�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ���?wqwq�?�T�H��?^�
�u��?7��XQ�?�@�Ե�?�������?333333�?      �?        �������?333333�?      �?                      �?#,�4�r�?�{a���?������?�}A_Ї?�������?������y?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?              �?|a���?	�=����?ZZZZZZ�?�������?              �?      �?      �?�s�9��?�c�1Ƹ?              �?�������?�?O��N���?;�;��?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?              �?      �?              �?      �?                      �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?              �?/�袋.�?F]t�E�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?              �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ"�hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         d                    �?���-�g�?�           ��@              S                    �?6�����?�            `v@              $                    �?2k��%�?�            �r@              #                 ���@p�eU}�?�            �i@                                  �?@���p��?�            `i@        ������������������������       �        /             R@                                   @M@�	a�$a�?X            ``@              	                    �?��:�-�?G            @Y@        ������������������������       �                     6@        
                          @[@pY���D�?8            �S@                                   �G@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                   @L@ �й���?4            @R@       ������������������������       �        /             P@                                   �L@�����H�?             "@                                 �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  `_@�������?             >@                                  �`@����X�?             @        ������������������������       �                     �?                                   �?r�q��?             @                                 @e@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                      
             �?���}<S�?             7@       ������������������������       �                     *@               "                    �?z�G�z�?             $@               !                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        %       H                    �?�W*��?B            @X@       &       +                    �D@L������?4            �S@        '       *                    �?�����H�?             "@        (       )                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ,       A                    �?B� ��?.            �Q@       -       2                    �?����0�?$             K@        .       1                    �?�8��8��?             (@        /       0                    s@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        3       6                    ]@և���X�?             E@        4       5                    �E@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        7       8                   @_@:ɨ��?            �@@        ������������������������       �                     @        9       @                   �d@PN��T'�?             ;@       :       ;                    @H@�<ݚ�?             2@        ������������������������       �                      @        <       =                    @N@      �?             0@       ������������������������       �        	             (@        >       ?                    �O@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        B       C                    �H@      �?
             0@        ������������������������       �                     @        D       E                   �n@$�q-�?	             *@       ������������������������       �                     $@        F       G                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        I       L                    �?X�<ݚ�?             2@       J       K                    T@      �?
             (@        ������������������������       �                     @        ������������������������       �                     "@        M       R                   �\@r�q��?             @       N       Q                    �?z�G�z�?             @       O       P                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        T       [                    �?t�6Z���?%            �K@        U       V                   �_@�q�q�?
             2@        ������������������������       �                      @        W       X                     L@���Q��?             $@        ������������������������       �                     @        Y       Z       
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        \       a                   �a@@-�_ .�?            �B@       ]       ^                   �c@      �?             @@       ������������������������       �                     <@        _       `                   �d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        b       c                   �U@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        e       �       	             �?�l�	jM�?�            �w@       f       �                    _@�[5]|x�?�            @v@        g       x                    �?      �?B             [@        h       s                    @M@      �?             @@       i       r                   pp@
;&����?             7@       j       m                   a@ҳ�wY;�?             1@        k       l                   �^@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        n       o                    �L@"pc�
�?             &@       ������������������������       �                      @        p       q                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       w                   �k@�����H�?             "@        u       v                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        y       ~                   �b@�=A�F�?-             S@       z       }                    �?�U�:��?"            �M@        {       |                    @H@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �I@               �                     D@j���� �?             1@        �       �       
             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @G@      �?             (@       ������������������������       �                      @        �       �                   �d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?T�AI-��?�             o@        �       �                    @G@ {��e�?D            �Z@        ������������������������       �                     @        �       �                   ph@tt���A�?C            �Y@        ������������������������       �                    �D@        �       �                    �?V��z4�?(             O@        �       �                    �?D�n�3�?             3@       �       �                   (s@"pc�
�?             &@       �       �                    n@ףp=
�?             $@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �N@      �?              @       �       �       
             �?      �?             @        ������������������������       �                     �?        �       �                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @H@�%^�?            �E@        ������������������������       �                     @        �       �                    �?z�G�z�?             D@        �       �                    �?ҳ�wY;�?             1@        �       �                   �^@և���X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @       �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �[@�z�G��?             $@        �       �                     J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���}<S�?             7@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                   `Z@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        �       �                    �?X�.�d�?W            �a@        �       �                    �?�חF�P�?             ?@       �       �                 ��� @z�G�z�?             9@       �       �                    �?�	j*D�?             *@       �       �                    �?X�<ݚ�?             "@        �       �                   @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@և���X�?             @        ������������������������       �                      @        �       �                   �`@���Q��?             @        ������������������������       �                      @        �       �                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `@�8��8��?             (@        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        D            �[@        �       �                   �^@�G�z��?             4@        ������������������������       �                     @        �       �                    �?d}h���?	             ,@       �       �                    @F@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  lk�w��?J��	.�?�*��o��?1��� ��?������?�+�Q���?(�J��"�?��VCӭ?�W�Δ�?xÏ���?      �?        T���0��?`�	)y��?0��<�]�?��be�F�?      �?        a~W��0�?�3���?�������?UUUUUU�?              �?      �?        ����Ǐ�?����?      �?        �q�q�?�q�q�?�������?�������?              �?      �?              �?        �������?�������?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?�������?�������?              �?      �?                      �?ӛ���7�?d!Y�B�?      �?        �������?�������?333333�?�������?              �?      �?              �?                      �?�Q�/�~�?_\����?h *�3�?1���M��?�q�q�?�q�q�?      �?      �?      �?                      �?              �?B�A��?|�W|�W�?�Kh/���?Lh/����?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?�q�q�?�q�q�?      �?                      �?N6�d�M�?e�M6�d�?              �?&���^B�?h/�����?9��8���?�q�q�?              �?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?r�q��?�q�q�?      �?      �?              �?      �?        UUUUUU�?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?��)A��?X���oX�?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?        �������?�������?      �?                      �?к����?S�n0E�?      �?      �?              �?      �?      �?      �?                      �?�������?�������?      �?                      �?�\AL� �?ڨ�l�w�?7��Mmj�?����d%�?      �?      �?      �?      �?�Mozӛ�?Y�B��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        /�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?6��P^C�?��k(��?�pR�屵?�A�I�?      �?      �?              �?      �?                      �?�������?ZZZZZZ�?�������?�������?              �?      �?              �?      �?      �?              �?      �?      �?                      �?�{��޻?�B!��?
�[���?~�	�[�?      �?        ��O ���?����?              �?�s�9��?2�c�1�?(������?l(�����?F]t�E�?/�袋.�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �}A_�?�}A_��?      �?        �������?�������?�������?�������?۶m۶m�?�$I�$I�?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        333333�?ffffff�?      �?      �?              �?      �?                      �?d!Y�B�?ӛ���7�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?�@�6�?�ۥ����?��RJ)��?�Zk����?�������?�������?;�;��?vb'vb'�?�q�q�?r�q��?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?�������?�������?              �?I�$I�$�?۶m۶m�?]t�E�?F]t�E�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���"hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKÅ�h��B�0         P                 ����?���-�g�?�           ��@              9                    �?�E����?�            �v@              6                    �?�uW��?�            `o@                                  P@ĴF���?�            �n@                                   �?�\��N��?             3@                                  @\@      �?              @              
                    �?�q�q�?             @              	                   p`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?���|���?             &@        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     @                                  @b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?               #                    �?`�F���?�            `l@                                  @L@ �.�?Ƞ?u            �f@       ������������������������       �        \            �b@                                   �L@ףp=
�?             >@                                   c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               "                    �N@@4և���?             <@              !       	             �?8�Z$���?             *@                                   @N@����X�?             @                                  �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        $       5       
             �?��k=.��?             �G@       %       0       	             �?8^s]e�?             =@       &       -                    �L@��S���?             .@       '       *                   `\@�q�q�?             "@        (       )                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        +       ,                   �c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        .       /                   f@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        1       2                    �?@4և���?             ,@        ������������������������       �                     �?        3       4                    d@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �        
             2@        7       8                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        :       ;                   ph@Rԅ5l�?F            @[@        ������������������������       �                     K@        <       O                    �?�b��[��?(            �K@       =       H                 ����?�+��<��?!            �E@       >       C                   �b@�<ݚ�?             ;@       ?       B                    @E@�C��2(�?             6@        @       A                     D@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     2@        D       E                   �d@z�G�z�?             @       ������������������������       �                     @        F       G       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J       
             �?     ��?             0@       ������������������������       �                     $@        K       L                    c@      �?             @        ������������������������       �                      @        M       N                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        Q       �       	             �?N�_����?�            `w@       R       {                    �?,�"���?�            @u@        S       z                   �s@Hg����?9            �V@       T       a                    �?H�U?B�?5            �T@        U       X                   �_@��
P��?            �A@        V       W                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        Y       `                   `f@��+7��?             7@       Z       ]                    �?��s����?             5@       [       \                    U@      �?             0@        ������������������������       �                      @        ������������������������       �        	             ,@        ^       _                 ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        b       y                   �c@��|�5��?            �G@       c       f                   �\@"pc�
�?             F@        d       e                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        g       x                 `ff�?�p ��?            �D@       h       m                    �?z�G�z�?             >@        i       j                   `Z@�q�q�?             @        ������������������������       �                     �?        k       l                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        n       q                 ����?�8��8��?             8@        o       p                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        r       w                    @N@P���Q�?             4@        s       t                 033�?ףp=
�?             $@        ������������������������       �                     @        u       v                   d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        |       �                    �? "��u�?�            @o@        }       ~                   �i@h㱪��?D            �[@        ������������������������       �                     C@               �                    @G@�X�<ݺ?-             R@        �       �                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�nkK�?+            @Q@       �       �                    �?�8���?#             M@       �       �                 ����? ��WV�?              J@        �       �                    �?r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     D@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   0k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    @N@���2���?W            �a@       �       �                    �?�Cc}h��?D             \@        �       �                   �w@��s����?             5@       �       �                   �U@�KM�]�?             3@        ������������������������       �                     �?        �       �                 `ff�?�X�<ݺ?             2@       ������������������������       �        	             *@        �       �                    �?z�G�z�?             @       �       �                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @M@$�q-�?6            �V@       �       �                   �r@����!p�?4             V@       �       �                   `_@xL��N�?+            �R@       ������������������������       �                    �E@        �       �                    �K@��a�n`�?             ?@       �       �                   �g@ 7���B�?             ;@        �       �                   �V@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             3@        �       �                    ^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ����?؇���X�?	             ,@        �       �                 ����?�q�q�?             @        ������������������������       �                     �?        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     <@        �       �                    @L@j���� �?             A@       �       �                    �?�q�q�?             8@        ������������������������       �                     @        �       �                   �d@�t����?
             1@       �       �                   �p@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B0  lk�w��?J��	.�?r�q��?�q�q�?���Q��?FA@s}�?E�JԮD�?ە�]�ڵ?y�5���?�5��P�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        F]t�E�?]t�E]�?              �?      �?      �?      �?        �������?�������?              �?      �?        �E�V�N�?E�����?wwwwww�?�?      �?        �������?�������?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?;�;��?;�;��?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?      �?              �?        g���Q��?br1���?|a���?	�=����?�������?�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?      �?        n۶m۶�?�$I�$I�?      �?        �؉�؉�?;�;��?      �?                      �?      �?        �������?�������?      �?                      �?�d	l�O�?���d	l�?              �?־a��?� O	��?w�qG�?w�qG��?�q�q�?9��8���?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?�������?�������?      �?              �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?      �?              �?      �?                      �?��/G��?�y4���?�������?�?��O��O�?�-؂-��?�v%jW��?�D�JԮ�?PuPu�?_�_��?UUUUUU�?UUUUUU�?      �?                      �?zӛ����?Y�B��?z��y���?�a�a�?      �?      �?              �?      �?        333333�?�������?              �?      �?                      �?x6�;��?br1���?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?��+Q��?Q��+Q�?�������?�������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?        �������?ffffff�?�������?�������?              �?�������?�������?              �?      �?                      �?              �?      �?              �?        ���Q��?�G�z�?��)A��?־a���?              �?�q�q�?��8��8�?UUUUUU�?UUUUUU�?      �?                      �?d!Y�B�?�Mozӛ�?a���{�?j��FX�?;�;��?O��N���?UUUUUU�?�������?              �?      �?                      �?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?�A�A�?�W|�W|�?I�$I�$�?�m۶m��?�a�a�?z��y���?(�����?�k(���?      �?        �q�q�?��8��8�?              �?�������?�������?      �?      �?              �?      �?                      �?      �?        ;�;��?�؉�؉�?]t�E�?/�袋.�?L�Ϻ��?>�S��?              �?�c�1Ƹ?�s�9��?h/�����?	�%����?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?ZZZZZZ�?UUUUUU�?�������?      �?        �������?�������?;�;��?;�;��?      �?                      �?      �?      �?      �?                      �?�������?�������?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�h�hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKɅ�h��B@2         d                    �?�ܲ�}��?�           ��@              Y       	             �?z0�R�W�?
           `y@              "                    �?�!�I�*�?�            �w@                                   �?nM`����?             G@                                  �?r֛w���?             ?@                                  �R@      �?             (@        ������������������������       �                     @               	                   @_@      �?              @        ������������������������       �                     @        
                           �?      �?             @                                 �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                  �`@�KM�]�?             3@                                  �?"pc�
�?             &@                                  �?�<ݚ�?             "@                                  �L@����X�?             @                                 h@      �?             @        ������������������������       �                     �?                                  �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @               !                   �a@���Q��?	             .@                                   �?ףp=
�?             $@                                  �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        #       N                    �?|�(8��?�            �t@       $       %                 ����?��/1��?�            t@        ������������������������       �        +            �P@        &       =       
             �?HVĮ���?�            �o@       '       <                    �R@P�S�L�?�            `j@       (       7                    �?@�S�1�?�             j@       )       *                   �V@F��}��?`            @b@        ������������������������       �                     �?        +       ,                 ����?�2c�$��?_             b@        ������������������������       �                     �?        -       4                   0j@ �q�q�?^             b@        .       /                   �h@�����H�?            �F@       ������������������������       �                    �C@        0       1                    ^@r�q��?             @        ������������������������       �                     @        2       3                 @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        5       6                 ����?`�LVXz�?A            �X@        ������������������������       �                     �?        ������������������������       �        @            �X@        8       ;                 ����? ������?,            �O@        9       :                    �?�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        ������������������������       �        !             G@        ������������������������       �                      @        >       I                    �?RB)��.�?            �E@       ?       H                    c@�c�Α�?             =@       @       E                   �m@�J�4�?             9@       A       B                   �b@���N8�?             5@       ������������������������       �        	             1@        C       D                     G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        F       G                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        J       M                 ����?@4և���?	             ,@        K       L                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        O       X                    �?�n_Y�K�?	             *@       P       Q                    �?X�<ݚ�?             "@        ������������������������       �                     �?        R       U                   �b@      �?              @        S       T                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        V       W                   Pp@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Z       [                   �^@R�}e�.�?             :@        ������������������������       �                     @        \       ]                   �\@��2(&�?             6@        ������������������������       �                     �?        ^       c                   pb@�����?             5@       _       `                 `ff�?P���Q�?
             4@       ������������������������       �                     1@        a       b                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        e       �                   �g@���O�`�?�            �t@       f       �                    �?P�4"7��?�            Pt@       g       p                    �?���T��?�            `q@        h       o                 033@P��BNֱ?1            �T@       i       j       
             �?��Y��]�?0            �T@       ������������������������       �                     L@        k       l                    �?$�q-�?             :@       ������������������������       �                     4@        m       n                     P@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        q       �                    �?�r����?v            `h@       r       �                   `@�KM�]�?i            `e@        s       �                    �?�z����?,            @P@        t       �                     L@�z�G��?             4@       u       �                    @�eP*L��?             &@       v       w                     D@�q�q�?             "@        ������������������������       �                     @        x                           p@���Q��?             @       y       ~                    �I@      �?             @       z       {                   �`@�q�q�?             @        ������������������������       �                     �?        |       }                    @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @33�?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   pj@�����H�?            �F@        ������������������������       �                     4@        �       �       
             �?z�G�z�?             9@       �       �                 ����?���y4F�?             3@       �       �                    @L@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @p@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pb@�8�l��?=            �Z@       �       �                    �?x�G�z�?.             T@        ������������������������       �                     1@        �       �                    �O@���N8�?#            �O@       �       �       	             �? _�@�Y�?              M@       �       �                    �?��?^�k�?            �A@        �       �                    �?�}�+r��?	             3@       ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �                     7@        �       �                 ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	             �?8�Z$���?             :@       �       �                    �L@������?	             .@       ������������������������       �                      @        �       �                    �?և���X�?             @       �       �                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?�q�q�?             8@       �       �                    �?���|���?             6@       �       �                 `ffֿ�E��ӭ�?	             2@        ������������������������       �                      @        �       �                 433�?     ��?             0@       �       �                   �`@@4և���?             ,@        �       �                    ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        �       �                 @33�?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?֭��F?�?            �G@        ������������������������       �                     *@        �       �                    �?��hJ,�?             A@       �       �                    @I@z�G�z�?             9@        �       �                    �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    `@��2(&�?             6@       ������������������������       �                     (@        �       �                   �b@�z�G��?             $@       �       �                 `ff�?      �?              @        �       �                    @K@z�G�z�?             @        ������������������������       �                     @        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ����u��?/�E��?"\E;�?}7��.1�?�ĩ�sK�?i�
��v�?zӛ����?C���,�?�B!��?���{��?      �?      �?              �?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        (�����?�k(���?F]t�E�?/�袋.�?�q�q�?9��8���?�$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?              �?333333�?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�!�c)�?�;�Ӛ�??q��z�?���R��?              �?
�B�P(�?_����z�?JQ/#��?`�
��T�?P���?�?G�<��?����?��Ǐ?�?      �?        �y�!���?cH�-�t�?      �?        UUUUUU�?�������?�q�q�?�q�q�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?[�R�֯�?�~�@��?      �?                      �?AA�?��}��}�?�?�?              �?      �?                      �?      �?        ���)k��?S֔5eM�?�{a���?5�rO#,�?{�G�z�?�z�G��?�a�a�?��y��y�?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?      �?        �$I�$I�?n۶m۶�?�������?�������?              �?      �?                      �?ى�؉��?;�;��?r�q��?�q�q�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?              �?'vb'vb�?�;�;�?              �?��.���?t�E]t�?              �?=��<���?�a�a�?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?���|�?���|��?��J�?�������?�"gXp��?��<}��?��FS���?���ˊ��?8��18�?������?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�?�k(���?(�����?[��Z���?�Z��Z��?ffffff�?333333�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?        �������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?              �?�q�q�?�q�q�?      �?                      �?�q�q�?�q�q�?      �?        �������?�������?6��P^C�?(������?      �?      �?      �?                      �?              �?�������?UUUUUU�?              �?      �?        �>����?�	�[��?�������?333333�?      �?        ��y��y�?�a�a�?#,�4�r�?�{a���?_�_��?�A�A�?�5��P�?(�����?      �?                      �?      �?              �?        333333�?�������?              �?      �?        ;�;��?;�;��?wwwwww�?�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?]t�E]�?F]t�E�?�q�q�?r�q��?              �?      �?      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?              �?      �?              �?        br1���?�F}g���?      �?        �������?KKKKKK�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        t�E]t�?��.���?              �?333333�?ffffff�?      �?      �?�������?�������?              �?      �?      �?      �?                      �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���RhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK酔h��B@:         j                 ����?({E�B��?�           ��@              +                    �?�V��?�            `w@                                   �?6�����?A            @[@                                   �J@և���X�?             5@                                  �?���Q��?
             .@        ������������������������       �                     @               
                    �F@���Q��?             $@               	       
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                      
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?h�V���?4             V@                                   �?���Q��?             @        ������������������������       �                      @                                  �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?               &       	             �?�+Ĺ+�?0            �T@                                  �O@      �?-             T@                                 �`@ ��ʻ��?$             Q@       ������������������������       �                     H@                                   �?P���Q�?             4@                                  d@@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     @               #                     P@�q�q�?	             (@               "                    �?      �?             @               !                    `@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        $       %                 ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        '       *                    �?�q�q�?             @       (       )                   0o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ,       Y                    �?����l�?�            �p@       -       0                   `X@��u}���?�            �m@        .       /                   �X@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        1       @                   @E@ ��Ou��?�            @m@        2       7                    �?�ՙ/�?             5@        3       4                    �?�C��2(�?             &@       ������������������������       �                     @        5       6                    `Q@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        8       9                   `[@�z�G��?             $@        ������������������������       �                      @        :       ?                    �?      �?              @       ;       >                 ����?؇���X�?             @        <       =                   Pa@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        A       R                     P@(�Y��E�?�            �j@       B       C                    �?�)f5��?�            �i@       ������������������������       �        q            �e@        D       I                    @F@�n`���?             ?@        E       H                   i@�q�q�?             "@        F       G       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        J       Q                   �g@��2(&�?             6@       K       L                    �?P���Q�?             4@       ������������������������       �                     &@        M       P                    �?�����H�?             "@        N       O                   d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        S       X                   @o@      �?              @       T       W       	             �?      �?             @       U       V                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Z       c                   �j@�q�q�?             ;@        [       b                 ����?և���X�?             @       \       ]                    a@      �?             @        ������������������������       �                     �?        ^       _                    �?�q�q�?             @        ������������������������       �                     �?        `       a                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        d       e                   `c@      �?             4@        ������������������������       �                     $@        f       g                    �?      �?             $@        ������������������������       �                      @        h       i                   Pd@      �?              @        ������������������������       �                     @        ������������������������       �                     @        k       �       
             �?R���Q�?�            �v@       l                           �?�o�����?�            �r@        m       p                    �?X�<ݚ�?             B@        n       o                 ���@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        q       ~       	             �?���Q��?             9@       r       w                   �q@����X�?             5@       s       v                    �?�8��8��?	             (@        t       u                     Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        x       }                 ����?X�<ݚ�?             "@       y       |                     L@r�q��?             @        z       {                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�K��G^�?�            @p@        �       �                    �?�����?             C@       �       �                    �?ҳ�wY;�?             A@       �       �                    �?"pc�
�?             6@       �       �                   pl@���y4F�?             3@        �       �                    �L@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �       �                   ``@�q�q�?             (@        ������������������������       �                     @        �       �                    d@�����H�?             "@       ������������������������       �                     @        �       �                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����?�            �k@        �       �                    �?r�q��?*             R@       �       �                    �?���5��?!            �L@        �       �                   �l@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�nkK�?             G@        �       �                    �M@�X�<ݺ?	             2@       ������������������������       �                     $@        �       �                   �`@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �c@h�����?             <@       ������������������������       �                     6@        �       �                   �r@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?	             .@       �       �                   �t@X�<ݚ�?             "@       �       �                    S@����X�?             @        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? "��u�?b            �b@        ������������������������       �                     8@        �       �                    �M@@4և���?Q            �_@       �       �                    c@ܷ��?��?9            �U@       �       �                   @\@�8��8��?7             U@        �       �                   �[@"pc�
�?             6@       �       �                    �?ףp=
�?             4@       ������������������������       �                     (@        �       �                   @^@      �?              @        ������������������������       �                     @        �       �                    b@���Q��?             @       �       �                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �h@Hn�.P��?+             O@        ������������������������       �                     8@        �       �                   @i@�˹�m��?             C@        ������������������������       �                      @        �       �                   �\@������?             B@        �       �                   p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �C@        �       �                   �d@     ��?+             P@        �       �                    �M@�IєX�?             1@       ������������������������       �                     (@        �       �                   @`@z�G�z�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�[�IJ�?            �G@       �       �                    �?�q�q�?            �C@        ������������������������       �                     @        �       �                    b@     ��?             @@       �       �                   ``@|��?���?             ;@       �       �                    �?�q�q�?             5@        ������������������������       �                     @        �       �                 ��� @j���� �?
             1@       �       �                   �b@      �?	             0@       �       �                   @_@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   i@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  Ac�Zb�?`yΨ�N�?�и[��?1�_�H1�?4R1�:#�?s�3R1��?۶m۶m�?�$I�$I�?333333�?�������?      �?        �������?333333�?333333�?�������?              �?      �?        �������?�������?      �?                      �?              �?/�袋.�?�袋.��?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���ˊ��?(፦ί�?      �?      �?�?�������?              �?�������?ffffff�?�$I�$I�?n۶m۶�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?���W��?үz�@�?�o��o��?�\�\�?      �?      �?              �?      �?        .��-���?�i�i�?�<��<��?�a�a�?]t�E�?F]t�E�?      �?        �������?�������?      �?                      �?333333�?ffffff�?      �?              �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�3����?��χӠ?��;�?��߁��?      �?        �9�s��?�c�1��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ��.���?t�E]t�?ffffff�?�������?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?      �?              �?      �?              �?      �?        �������?�������?�n0E>��?S�n0E�?r�q��?�q�q�?]t�E�?F]t�E�?      �?                      �?�������?333333�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?r�q��?�q�q�?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?        �?�?�??�?��?^Cy�5�?Q^Cy��?�������?�������?F]t�E�?/�袋.�?(������?6��P^C�?�$I�$I�?۶m۶m�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?v�)�Y7�?�Ϻ���?UUUUUU�?�������?��Gp�?�}��?]t�E�?t�E]t�?              �?      �?        d!Y�B�?�Mozӛ�?�q�q�?��8��8�?              �?      �?      �?      �?      �?      �?                      �?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�q�q�?r�q��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?�������?      �?                      �?���Q��?�G�z�?              �?�$I�$I�?n۶m۶�?a���{�?��=���?UUUUUU�?UUUUUU�?F]t�E�?/�袋.�?�������?�������?              �?      �?      �?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �c�1ƨ?t�9�s�?              �?^Cy�5�?��P^Cy�?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�?�?              �?�������?�������?              �?      �?      �?      �?                      �?���
b�?m�w6�;�?UUUUUU�?UUUUUU�?      �?              �?      �?{	�%���?	�%����?UUUUUU�?UUUUUU�?      �?        �������?ZZZZZZ�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5\hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         Z                    �?�3u���?�           ��@                                  �?�b��-8�?�            �w@                      	             �?"pc�
�?%            �K@                                  �?f1r��g�?#            �J@                                   K@>a�����?"            �I@                                   �F@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        	                          �x@P���Q�?             D@       
                          �r@ ���J��?            �C@       ������������������������       �                     A@                                  �c@z�G�z�?             @        ������������������������       �                      @                                  �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               )                    �?@�0�!��?�            0t@              (                 ���@��$xtW�?�            �j@                                  @L@�n����?�            �i@                                 @g@PA��ڡ?i             e@                                 @[@�E��La�?h            �d@                      
             �?�����H�?             "@       ������������������������       �                     @                                  `m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        c            �c@        ������������������������       �                      @                '                    �M@�KM�]�?             C@        !       $                   �?����X�?             ,@        "       #                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        %       &                 ����?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     @        *       G                   �?���Q��?C            �[@       +       B                    �M@<ݚ)�?,             R@       ,       1                   �b@�z�6�?&             O@       -       .                    �?��?^�k�?            �A@       ������������������������       �                     8@        /       0                    @D@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        2       ?                   ``@X�<ݚ�?             ;@       3       :                    �?     ��?
             0@        4       9                    �?      �?              @       5       8                 ����?և���X�?             @       6       7                    e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ;       <                    @I@      �?              @       ������������������������       �                     @        =       >                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @       A                   �b@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        C       D                    �N@ףp=
�?             $@        ������������������������       �                     @        E       F                   Pd@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        H       M                 ����?D�n�3�?             C@        I       L                    �?z�G�z�?             $@       J       K                   `X@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        N       U                    �?      �?             <@        O       T                    �?     ��?             0@       P       S                 `ff@d}h���?             ,@       Q       R                   �k@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        V       Y                   �Y@�8��8��?	             (@        W       X                     M@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        [       �       
             �?�Mõ��?�            @v@       \       q                    �? U��?�            �q@        ]       p                    �?��V#�?            �E@       ^       o                     Q@؀�:M�?            �B@       _       `                   @[@^������?            �A@        ������������������������       �                     @        a       j                   �a@���Q��?             >@       b       c                 833�?     ��?             0@        ������������������������       �                      @        d       e                    �C@d}h���?
             ,@        ������������������������       �                      @        f       g                    @K@�8��8��?	             (@       ������������������������       �                     @        h       i                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        k       n                   `c@@4և���?	             ,@       l       m                     K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        r       �                   �f@X{����?�             n@       s       t                   �f@�e)���?�            �m@        ������������������������       �        /             Q@        u       �                 ����?��C[���?g             e@        v       �       	             �?h��Q(�?(            �P@       w       |                    �?\-��p�?#             M@        x       {                    �?�q�q�?             @       y       z                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        }       �                    �?X�;�^o�?             �K@       ~       �                   xp@��r._�?            �D@              �                   �o@�q�q�?             8@       �       �                    �?��s����?             5@       �       �                    �?���y4F�?             3@        �       �                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@�0�!��?
             1@       �       �                 ����?�8��8��?             (@       ������������������������       �                     @        �       �                   �j@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                    @I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             1@        ������������������������       �        	             ,@        �       �                   �_@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@@��j$޷??            �Y@       �       �                 ����?����?�?5            �V@        �       �                    �?@4և���?             <@       �       �                 033�?�����H�?             2@       ������������������������       �                     (@        �       �                     L@�q�q�?             @        ������������������������       �                     @        �       �                    �N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        %             O@        �       �                   �\@      �?
             (@        ������������������������       �                      @        �       �                    `@ףp=
�?             $@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����?b�2�tk�?/             R@        �       �                    �?�t����?             1@       �       �                    �?      �?             0@        �       �                    @F@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �F@\�����?"            �K@        ������������������������       �                     $@        �       �                   Pn@�L�lRT�?            �F@       �       �                    �?`՟�G��?             ?@        �       �                   �b@      �?              @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   P`@8����?             7@        �       �                    �?      �?              @       �       �                   �?և���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       �       �                     M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�r����?
             .@        �       �                    ]@      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                      @        �       �                   �Y@z�G�z�?             @       �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����?؇���X�?             ,@        �       �                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  k�w죻�?��	."�?�u]�u]�?QEQE�?F]t�E�?/�袋.�?�x+�R�?�!5�x+�?�?�������?t�E]t�?]t�E�?              �?      �?        �������?ffffff�?�A�A�?��-��-�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ZZZZZZ�?�������?����?��n�?�?�<����?j6��bP�?��s�n�?&�q-�?��4���?J����x?�q�q�?�q�q�?      �?              �?      �?      �?                      �?      �?                      �?�k(���?(�����?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?      �?              �?      �?              �?                      �?333333�?�������?��8��8�?�8��8��?J)��RJ�?�Zk����?_�_��?�A�A�?      �?        ]t�E�?F]t�E�?              �?      �?        r�q��?�q�q�?      �?      �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?]t�E�?F]t�E�?      �?                      �?�������?�������?              �?�������?�������?              �?      �?        (������?l(�����?�������?�������?�$I�$I�?�m۶m��?              �?      �?                      �?      �?      �?      �?      �?I�$I�$�?۶m۶m�?;�;��?;�;��?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?                      �?v�{��^�?#�E(�?�6��?�z2~���?6eMYS��?eMYS֔�?v�)�Y7�?E>�S��?_�_��?uPuP�?              �?�������?333333�?      �?      �?              �?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?�$I�$I�?n۶m۶�?UUUUUU�?�������?      �?                      �?              �?      �?                      �?ynyn�?�0��0��?�Ӭ����?�e��Ao�?              �?�B���Ǽ?�wɃg�?z�rv��?�Wc"=P�?�{a���?a����?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?J��yJ�?�־a��?ە�]���?�ڕ�]��?�������?�������?�a�a�?z��y���?(������?6��P^C�?      �?      �?              �?      �?        �������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �?nnnnnn�?l�l��?��I��I�?�$I�$I�?n۶m۶�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        9��8���?�8��8��?�?<<<<<<�?      �?      �?UUUUUU�?�������?      �?                      �?              �?      �?        A��)A�?߰�k��?      �?        l�l��?�I��I��?�s�9��?�1�c��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        8��Moz�?d!Y�B�?      �?      �?�$I�$I�?۶m۶m�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �?�������?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?              �?      �?                      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�Q&hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKυ�h��B�3         �                    �?�/�$�y�?�           ��@              K                    �?9h��S�?           @{@              >                    �?Riv����?�             r@                                  �?8��d�?�             o@                               033@����a�?v            `f@                                  �?�;Y�&��?u            @f@        ������������������������       �        '            �M@                                  @[@��u}���?N            �]@        	       
       	             �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @                                  �p@ \sF��?K            @\@                                  @L@@uvI��?A            �X@       ������������������������       �        5             T@                                  `a@�X�<ݺ?             2@       ������������������������       �                     $@                                   �?      �?              @        ������������������������       �                     @                                pff�?z�G�z�?             @                                 0b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                      
             �?������?
             .@                                  �?���Q��?             $@                                 �q@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                )                    �?&�a2o��?,            @Q@        !       $                   `\@$��m��?             :@        "       #                    �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        %       &                    r@�r����?             .@       ������������������������       �        	             (@        '       (                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        *       ;                    `P@�T|n�q�?            �E@       +       0                    �E@�ݜ�?            �C@        ,       /                   @b@�q�q�?             (@       -       .                    �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        1       2                    �I@ 7���B�?             ;@        ������������������������       �                     *@        3       :                   @`@@4և���?	             ,@        4       5                    �?z�G�z�?             @        ������������������������       �                      @        6       7                   Ph@�q�q�?             @        ������������������������       �                     �?        8       9                    n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        <       =                   @[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ?       J                 ����?��6���?             E@       @       A                    @E@�������?             >@        ������������������������       �                     @        B       I                   �_@HP�s��?             9@        C       D                    �z�G�z�?             $@        ������������������������       �                     �?        E       F                    �?�����H�?             "@        ������������������������       �                     @        G       H                    ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@        ������������������������       �                     (@        L       w                    �?`K�����?X            @b@        M       X                   �a@և���X�?+            �O@        N       S                   pm@���y4F�?             3@        O       R       	             �?      �?             @       P       Q                   `j@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        T       W                    Y@$�q-�?             *@        U       V                    �M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Y       ^                    �?d�
��?             F@        Z       ]                   �g@ףp=
�?	             $@        [       \                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        _       n       	             �?j���� �?             A@       `       e                    �? �o_��?             9@       a       d                   m@z�G�z�?
             .@       b       c                    @N@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        f       g                    ]@���Q��?             $@        ������������������������       �                     @        h       i                   �b@և���X�?             @        ������������������������       �                      @        j       k                   �`@z�G�z�?             @        ������������������������       �                     @        l       m                   @c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        o       r                    �?�<ݚ�?             "@        p       q                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       v                   �^@r�q��?             @        t       u                     D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        x                           �?��Lɿ��?-            �T@        y       z                 ����?��
ц��?             *@        ������������������������       �                     @        {       ~                    �N@�<ݚ�?             "@       |       }                    @L@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 033�?��?^�k�?'            �Q@       �       �                    �?@-�_ .�?            �B@       ������������������������       �                     >@        �       �                   o@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �@@        �       �                    �?�`
\b�?�            �r@        �       �                    @K@���3�E�?#             J@        �       �                    �?�ՙ/�?             5@       �       �                    V@�θ�?	             *@        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �k@      �?              @        �       �       	             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?`Jj��?             ?@       ������������������������       �                     :@        �       �                   �b@���Q��?             @       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?������?�            �n@       �       �                    �?���Hx�?�             k@        �       �                    �?4�2%ޑ�?            �A@        �       �                   �b@�<ݚ�?             "@        ������������������������       �                     @        �       �                     M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �? ��WV�?             :@        �       �                    @M@z�G�z�?             @       �       �                    f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             5@        �       �                    `@�����?m            �f@       �       �                 ����?؀���˲?P            ``@        �       �                    Z@�U�:��?!            �M@        ������������������������       �        	             7@        �       �                    �?4?,R��?             B@        �       �                    �M@���Q��?             @       �       �                    ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    \@`Jj��?             ?@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     7@        ������������������������       �        /             R@        �       �                 ����?�J�4�?             I@        �       �                    �?�t����?             1@        �       �                   pl@      �?             $@        �       �                     L@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @b@�C��2(�?            �@@       �       �                 ����? ��WV�?             :@        �       �                   0j@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             4@        �       �                 `ff�?����X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    W@ףp=
�?             >@        ������������������������       �                     �?        �       �                     R@ 	��p�?             =@       ������������������������       �                     ;@        ������������������������       �                      @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B�  L�f���?Z�L��?��ش��?	l�O���?>�����?	�=����?��RJ)��?�Zk��ֺ?����X6�?�Fu��?�0�9�a�?��g<�?      �?        �o��o��?�\�\�?UUUUUU�?UUUUUU�?              �?      �?        [X驅��?Vzja���?�Cc}h��?9/���?      �?        ��8��8�?�q�q�?      �?              �?      �?      �?        �������?�������?      �?      �?              �?      �?              �?        wwwwww�?�?333333�?�������?      �?      �?              �?      �?                      �?      �?                      �?��Q�g��?ہ�v`��?�N��N��?vb'vb'�?F]t�E�?]t�E]�?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?���)k��?6eMYS��?\��[���?�i�i�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?	�%����?h/�����?      �?        n۶m۶�?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?      �?      �?                      �?b�a��?=��<���?�������?�������?              �?q=
ףp�?{�G�z�?�������?�������?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?����Ǐ�?���?۶m۶m�?�$I�$I�?(������?6��P^C�?      �?      �?      �?      �?              �?      �?              �?        ;�;��?�؉�؉�?�������?�������?      �?                      �?              �?�袋.��?�.�袋�?�������?�������?      �?      �?      �?                      �?      �?        ZZZZZZ�?�������?�Q����?
ףp=
�?�������?�������?      �?      �?              �?      �?                      �?�������?333333�?              �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?              �?      �?              �?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        rY1P»?�������?�;�;�?�؉�؉�?              �?9��8���?�q�q�?333333�?�������?      �?                      �?      �?        �A�A�?_�_��?к����?S�n0E�?              �?�$I�$I�?�m۶m��?      �?                      �?              �?i���m��?&����?b'vb'v�?O��N���?�<��<��?�a�a�?ى�؉��?�؉�؉�?              �?      �?              �?      �?333333�?�������?              �?      �?                      �?�B!��?���{��?              �?�������?333333�?      �?      �?      �?                      �?      �?        ������?�|����?9��8��?9��8���?�A�A�?�������?9��8���?�q�q�?      �?        333333�?�������?      �?                      �?;�;��?O��N���?�������?�������?      �?      �?              �?      �?                      �?              �?�jc�?]��ҟ��?�i��?h�T��?�pR�屵?�A�I�?              �?r�q��?�8��8��?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �B!��?���{��?      �?      �?              �?      �?                      �?              �?{�G�z�?�z�G��?�������?�������?      �?      �?�m۶m��?�$I�$I�?      �?                      �?              �?              �?F]t�E�?]t�E�?;�;��?O��N���?UUUUUU�?�������?      �?                      �?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        �{a���?������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ&N�hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKㅔh��B�8         �                    �?p�Vv���?�           ��@              I                   �a@�Y����?           �z@              2                 pff�?�luL3�?�            Ps@               +                    �N@����>4�?O             \@              "                    �?ڤ���?9            @T@                                  �?r�z-��?%            �J@                                  �v@"pc�
�?             &@                                  �?ףp=
�?             $@        	       
       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                   �?d}h���?             E@                     	             �?���}<S�?             7@       ������������������������       �                     3@                                  `Y@      �?             @        ������������������������       �                     �?                                  �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �g@p�ݯ��?             3@        ������������������������       �                     @                                   �?��
ц��?	             *@        ������������������������       �                     �?                                   �?�q�q�?             (@        ������������������������       �                     @                                  �\@X�<ݚ�?             "@        ������������������������       �                      @                                  �j@����X�?             @        ������������������������       �                     �?                !                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        #       $                 ����?@4և���?             <@       ������������������������       �                     5@        %       *                    �?����X�?             @       &       )                    �?���Q��?             @       '       (                    n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ,       /                   P`@`Jj��?             ?@       -       .                    �R@XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        0       1                     Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       B                 pff�?��I�~R�?n            �h@        4       A                   �j@     ��?&             P@        5       6                    �?�S����?             C@        ������������������������       �                     @        7       >                   �c@�IєX�?             A@       8       9                    �?      �?             @@       ������������������������       �                     6@        :       ;                     O@ףp=
�?             $@        ������������������������       �                      @        <       =                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ?       @                 pff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        C       H                    �?pJQg���?H            �`@        D       E                    @P@ףp=
�?             >@       ������������������������       �                     7@        F       G                     Q@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        9            �Y@        J       �                    �?�n\�GZ�?I            �]@       K       |                   �q@X�����?7             V@       L       u       	             �?L�];�?-            �Q@       M       t                    �O@D7�J��?#            �K@       N       e       
             �?և���X�?             �H@       O       X                   Ph@¦	^_�?             ?@        P       W                    �?�z�G��?             $@       Q       V                   `e@�<ݚ�?             "@       R       S                    �?      �?              @        ������������������������       �                     @        T       U                 ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                   �_@�����?             5@        ������������������������       �                     &@        [       ^                    �?z�G�z�?             $@        \       ]                   Pp@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                 033�?      �?              @        ������������������������       �                     @        a       d                   �a@z�G�z�?             @        b       c                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        f       s                    �?�q�q�?             2@       g       l                   Ph@      �?
             (@        h       k                   �`@      �?             @       i       j                   �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        m       n                     G@      �?              @        ������������������������       �                     @        o       r                    �?���Q��?             @       p       q                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        v       y                    �K@      �?
             0@       w       x                    �?@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        z       {                 hff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        }       �                    �E@�t����?
             1@        ~                           �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        �       �                 033@��a�n`�?             ?@       �       �                    @L@h�����?             <@        �       �                   �m@؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        �       �                   `e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @E@��S����?�             s@        �       �                 833�?     ��?             @@        �       �                    a@�eP*L��?             &@       �       �                    �?�q�q�?             "@       �       �                    �P@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �M@؇���X�?             5@       ������������������������       �                     1@        �       �                   `V@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?d/�@7�?�             q@       �       �                    �?������?h             c@       �       �                   �b@��d��?U            �_@       �       �                    @ ��(��?L            @\@       �       �       
             �?��#:���?J            �[@       �       �                   �b@�����D�?*            @P@       �       �                   Pa@�(\����?             D@       ������������������������       �                     5@        �       �                   �o@�}�+r��?             3@       ������������������������       �                     0@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   @c@� �	��?             9@        ������������������������       �                      @        �       �                    k@�û��|�?             7@        �       �                   pe@�z�G��?             $@       �       �                    �?؇���X�?             @       �       �                   pj@r�q��?             @       �       �                     E@�q�q�?             @        ������������������������       �                     �?        �       �                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �n@8�Z$���?	             *@       ������������������������       �                     @        �       �                   `o@�q�q�?             @        ������������������������       �                     �?        �       �                   �d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�����H�?             �F@       �       �                   @[@      �?             D@        �       �                   @Z@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�8��8��?             B@       �       �                   Pc@��2(&�?             6@       ������������������������       �        
             &@        �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �                    a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             *@        �       �                    �?�5��?             ;@       �       �                    �?z�G�z�?
             .@       �       �                 033�?�z�G��?             $@       �       �                   �e@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�q�q�?	             (@       �       �                    �?      �?              @        ������������������������       �                     �?        �       �                 033�?և���X�?             @       �       �                    �?      �?             @       �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        C            @^@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  w
��,@�?�z�����?&�;u-�?���4>�?NZ�Ϯ�?�+&��?I�$I�$�?n۶m۶�?X�<ݚ�?����H�?�琚`��?����!�?/�袋.�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?۶m۶m�?I�$I�$�?d!Y�B�?ӛ���7�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        Cy�5��?^Cy�5�?              �?�;�;�?�؉�؉�?              �?�������?�������?      �?        �q�q�?r�q��?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?�$I�$I�?n۶m۶�?              �?�$I�$I�?�m۶m��?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�B!��?���{��?�{a���?GX�i���?              �?      �?              �?      �?              �?      �?        \e
�d�?�Y���?      �?      �?^Cy�5�?(������?      �?        �?�?      �?      �?              �?�������?�������?              �?      �?      �?      �?                      �?      �?      �?              �?      �?                      �?�qA��?s���7G�?�������?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?              �?�O��O��?4X�3X��?F]t�E�?]t�E]�?SO�o�z�?Zas �
�?k߰�k�?J��yJ�?۶m۶m�?�$I�$I�?�RJ)���?��Zk���?ffffff�?333333�?9��8���?�q�q�?      �?      �?      �?              �?      �?              �?      �?                      �?              �?�a�a�?=��<���?              �?�������?�������?      �?      �?              �?      �?              �?      �?              �?�������?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?        �������?333333�?      �?      �?      �?                      �?              �?      �?              �?              �?      �?n۶m۶�?�$I�$I�?      �?                      �?      �?      �?      �?                      �?�?<<<<<<�?      �?      �?      �?                      �?              �?�c�1Ƹ?�s�9��?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?*�)��?Y�X��?      �?      �?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �ǭ��?��;�H��?xxxxxx�?�?��뺮��?EQEQ�?ja��V�?Vzja���?k߰��?�S�<%��?z�z��?z�z��?333333�?�������?      �?        �5��P�?(�����?      �?        UUUUUU�?UUUUUU�?      �?                      �?�Q����?)\���(�?              �?8��Moz�?��,d!�?333333�?ffffff�?�$I�$I�?۶m۶m�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?��.���?t�E]t�?      �?        F]t�E�?t�E]t�?      �?              �?      �?      �?                      �?      �?              �?                      �?      �?        /�����?h/�����?�������?�������?333333�?ffffff�?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��8hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B@/         V                    �?�3u���?�           ��@              I       	             �?>���Rp�?�            �w@              *                    �?�,�?2�?�            @o@              )                 ���@�j��e�?p            �f@                               ���ٿ��hJ,�?k            @e@        ������������������������       �                     @                                  @E@��(�#H�?i            �d@               	                     F@b�2�tk�?             2@        ������������������������       �                     @        
                          `_@��
ц��?	             *@                                  �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                  �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                  c@�m�&��?]            �b@                                   �?�\=lf�?,            �P@       ������������������������       �        (             O@                                   �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?               (       
             �?,���i�?1            �T@               '                    �?     ��?             @@                                 �c@��}*_��?             ;@        ������������������������       �                     @               &                    �?��+7��?             7@              %                   `m@���!pc�?             6@              $                     I@      �?             (@              #                    a@      �?              @              "                    �?؇���X�?             @               !                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     I@        ������������������������       �                     &@        +       .                    �?�G�5��?-            @Q@        ,       -                    �?�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        /       H                   Pd@�S����?&            �L@       0       9                    �?X�;�^o�?$            �K@       1       2                    �?(;L]n�?             >@        ������������������������       �                     �?        3       4                   �r@XB���?             =@       ������������������������       �                     9@        5       6                    �?      �?             @        ������������������������       �                     �?        7       8                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        :       C                    b@�+e�X�?             9@       ;       B                    �?R���Q�?             4@       <       A                 `ff�?�θ�?	             *@       =       >                   �^@�C��2(�?             &@       ������������������������       �                      @        ?       @                   �o@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        D       E                   �b@���Q��?             @        ������������������������       �                      @        F       G                   �e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        J       O                    I@�U���?L            �_@        K       L                    �?z�G�z�?             @        ������������������������       �                      @        M       N                   a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        P       Q                   �?��v$���?H            �^@       ������������������������       �        @             [@        R       U                   �_@؇���X�?             ,@        S       T                 pff�?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        W       n                    �?"oI���?�            Pv@        X       k                   �r@J�8���?(             M@       Y       b                    �?D^��#��?            �D@       Z       a                    �?z�G�z�?             4@       [       `                    �?�	j*D�?	             *@       \       ]                    [@      �?             (@        ������������������������       �                      @        ^       _                   �b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        c       j                   �a@؇���X�?             5@        d       e                   �\@���!pc�?             &@        ������������������������       �                     @        f       i                    k@      �?             @        g       h                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        l       m                   �c@�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        o       �                   `_@T�(�qu�?�            �r@        p       �                    �?\��<�|�?;            �W@        q       �       	             �?�\��N��?             C@       r       s                 @33�?�n_Y�K�?             :@        ������������������������       �                     $@        t                           �?      �?
             0@       u       |                    �?�eP*L��?             &@       v       w                    ]@      �?             @        ������������������������       �                      @        x       y                    �?      �?             @        ������������������������       �                      @        z       {                   m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        }       ~                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @I@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �^@�q�q�?             (@       �       �                    �?���Q��?             $@       �       �                    @H@z�G�z�?             @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?x�}b~|�?%            �L@       �       �                 ����?X�EQ]N�?            �E@        ������������������������       �                     3@        �       �                    �?�q�q�?             8@        �       �                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?      �?	             0@        �       �                    Y@�q�q�?             @        ������������������������       �                     �?        �       �                    �B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        
             ,@        �       �                    �?�IєX�?�            �i@        �       �                    �?�8��8N�?>             X@        �       �                    �?�+e�X�?             9@       �       �                    �I@z�G�z�?             4@        ������������������������       �                      @        �       �                    @�����H�?             2@       �       �                   �T@�IєX�?             1@        �       �                   �e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     �?        �       �                   �c@���Q��?             @       �       �                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   `X@ ��PUp�?)            �Q@        �       �                   �g@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        %            �O@        �       �       	             �?X'"7��?F             [@       �       �                    �?��s�n�?B             Z@       �       �                 ����?�ӖF2��?+            �Q@        �       �                 ����?������?
             1@       ������������������������       �                     *@        ������������������������       �                     @        �       �                   P`@@3����?!             K@        �       �                    �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                    �E@        ������������������������       �                    �@@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  k�w죻�?��	."�?�i��F�?GX�i���?#��~j��?�I+��?Ǉ 妢�?��}kdu�?KKKKKK�?�������?              �?�}�z���?3	v���?9��8���?�8��8��?              �?�;�;�?�؉�؉�?�$I�$I�?�m۶m��?      �?                      �?�������?UUUUUU�?      �?                      �?�?��8��?p�j:�?"=P9���?g��1��?      �?        �������?�������?      �?                      �?�����?8��18�?      �?      �?_B{	�%�?B{	�%��?              �?zӛ����?Y�B��?F]t�E�?t�E]t�?      �?      �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?              �?      �?              �?              �?              �?                      �?�%~F��?��v`��?UUUUUU�?UUUUUU�?      �?                      �?^Cy�5�?(������?J��yJ�?�־a��?�?�������?              �?�{a���?GX�i���?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ���Q��?R���Q�?333333�?333333�?�؉�؉�?ى�؉��?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ����|>�?��`0�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        .�u�y�?;ڼOqɐ?      �?        ۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?              �?      �?              �?        �J��J��?[�[��?|a���?�rO#,��?�]�ڕ��?,Q��+�?�������?�������?vb'vb'�?;�;��?      �?      �?              �?�������?�������?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?t�E]t�?F]t�E�?              �?      �?      �?      �?      �?              �?      �?              �?                      �?�?�?              �?      �?        V�)p��?u���A�?��%N��?��v�@�?�5��P�?y�5���?ى�؉��?;�;��?              �?      �?      �?t�E]t�?]t�E�?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?333333�?�������?      �?                      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?333333�?�������?�������?�������?      �?      �?      �?                      �?              �?      �?              �?        Lg1��t�?�YLg1�?qG�wĽ?w�qG�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?                      �?              �?�?�?�������?�������?���Q��?R���Q�?�������?�������?      �?        �q�q�?�q�q�?�?�?      �?      �?              �?      �?                      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?��V،?��ۥ���?      �?      �?              �?      �?                      �?B{	�%��?Lh/����?ى�؉��?b'vb'v�?�@�6�?�K=��?�?xxxxxx�?              �?      �?        h/�����?���Kh�?F]t�E�?]t�E�?      �?                      �?              �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�b�hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B@0         l                    �?�+	G�?�           ��@              S                    �?b���ނ�?           �z@                                 �Z@DѱS�7�?�            �t@                                   �?�t����?	             1@                                 �q@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     @        	       J                 033�?��z�H�?�            �s@       
       '                    �?|�����?�            �q@                                   �?f�<�>��?%            �M@                                ����?�>����?             ;@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �b@`2U0*��?             9@       ������������������������       �                     8@        ������������������������       �                     �?                                   �?     ��?             @@        ������������������������       �                      @               "                 ����?�q�q�?             >@                     	             �?"pc�
�?             6@                                  d@�KM�]�?             3@       ������������������������       �        	             &@                                ����?      �?              @                                  �?���Q��?             @        ������������������������       �                     �?                                  pd@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                !                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #       &       
             �?      �?              @       $       %                   Pp@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        (       A                    �?�&xw���?�            @l@       )       >                     R@��4+̰�?~            @h@       *       7                   �f@��8����?|             h@       +       0                   @[@�x�V�?v             g@        ,       /                    @I@�r����?             .@       -       .       
             �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        1       6                    �E@@c����?n            @e@        2       5                    _@@��8��?              H@        3       4                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     G@        ������������������������       �        N            �^@        8       9                    �?����X�?             @        ������������������������       �                     @        :       ;                   �g@      �?             @        ������������������������       �                     �?        <       =       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ?       @                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        B       I       	             �?     ��?             @@       C       D                    �?�q�q�?             8@        ������������������������       �                     "@        E       F                    @F@��S���?             .@        ������������������������       �                     @        G       H                    �M@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        K       R                    �?\-��p�?             =@        L       M                    �?      �?              @        ������������������������       �                     @        N       O                     P@z�G�z�?             @        ������������������������       �                      @        P       Q                   Pe@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        T       _                    �?�?�Ʋ(�?7            @W@        U       \       
             �?��
ц��?            �C@       V       [                 `ff�?      �?             @@       W       X                    ����N8�?
             5@        ������������������������       �                      @        Y       Z                    @E@�S����?	             3@        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     &@        ]       ^                   @V@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        `       a                     K@�>����?!             K@        ������������������������       �                     1@        b       k                    �?������?            �B@        c       h                   �b@������?	             1@       d       e                 ����?�8��8��?             (@       ������������������������       �                      @        f       g                   8p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        i       j                    e@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     4@        m       �                    �?��ѝ-�?�            `s@        n       �                   pa@l��[B��?$             M@       o       z                 ����?�Gi����?            �B@       p       y                    `P@p�ݯ��?             3@       q       x                     N@      �?             ,@       r       u                    �?�z�G��?             $@       s       t                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        v       w                   @^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        {       ~                   0a@r�q��?             2@       |       }                    �?@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?               �                   �l@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�ՙ/�?             5@        ������������������������       �                      @        �       �                    �?�n_Y�K�?             *@       �       �                   `c@      �?              @        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?$Q�q�?�            �o@       �       �                    \@ 7���B�?�             k@        �       �                   ``@��S�ۿ?.            �R@        �       �                    �?z�G�z�?             9@       �       �                   �[@���N8�?             5@       �       �                    @L@z�G�z�?             4@       �       �                    �I@@4և���?             ,@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?      �?             @       �       �                    �L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     I@        �       �                    Z@`Ql�R�?Z            �a@        �       �                   �a@      �?             @        ������������������������       �                     �?        �       �                    �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��[����?W             a@       �       �                 ����?@�n���?F            �Y@        �       �                    @G@������?             B@        �       �                    �?@4և���?	             ,@        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     6@        ������������������������       �        ,            �P@        ������������������������       �                     A@        �       �                 ����?�<ݚ�?             B@        �       �                    �D@�eP*L��?             &@        ������������������������       �                      @        �       �                    h@�q�q�?             "@        �       �                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `ff�?HP�s��?             9@       ������������������������       �                     7@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B  ��C�l�?z?+^���?��sH�?�9�&o�?9b�N���?wr�Ɲ�?�������?�������?;�;��?�؉�؉�?              �?      �?              �?        �a��x��?�x�YF�?��Q)z��?�	�Z��?�"h8���?��/���?�Kh/��?h/�����?      �?      �?      �?                      �?���Q��?{�G�z�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?F]t�E�?/�袋.�?(�����?�k(���?              �?      �?      �?�������?333333�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?333333�?�������?              �?      �?              �?        v��\�(�?�8�1�s�?_\����? tT����?�����*�?�������?��5!({�?�	A����?�������?�?�m۶m��?�$I�$I�?      �?                      �?      �?        �������?x?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?      �?�������?�������?      �?        �?�������?              �?F]t�E�?t�E]t�?      �?                      �?      �?        �{a���?a����?      �?      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?4�DM4�?f�]v�e�?�;�;�?�؉�؉�?      �?      �?�a�a�?��y��y�?              �?(������?^Cy�5�?              �?      �?                      �?�m۶m��?�$I�$I�?              �?      �?        h/�����?�Kh/��?              �?к����?��g�`��?�?xxxxxx�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?333333�?�������?      �?                      �?              �?+�"�*�?u;T�Cu�?GX�i���?���=��?#�u�)��?o0E>��?^Cy�5�?Cy�5��?      �?      �?ffffff�?333333�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?�������?�$I�$I�?n۶m۶�?              �?      �?              �?      �?      �?                      �?�<��<��?�a�a�?      �?        ى�؉��?;�;��?      �?      �?      �?      �?              �?      �?                      �?�������?�������?      �?                      �?AA�?~��}���?h/�����?	�%����?�?�������?�������?�������?��y��y�?�a�a�?�������?�������?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?                      �?      �?                      �?              �?W�+�ɕ?}g���Q�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ������}?�8R4��?��,�?\mMw��?�q�q�?�q�q�?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?              �?              �?              �?�q�q�?9��8���?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        {�G�z�?q=
ףp�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��bhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�6         x                    �?.��X~��?�           ��@                                 �\@�jTM��?�            �v@               
                 ����?���?            �D@                                   �?�z�G��?             $@                                  �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               	                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   @P@��a�n`�?             ?@                                  �?h�����?             <@       ������������������������       �        
             1@                                   �J@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                                   �?�q�q�?             @        ������������������������       �                     �?                                   �R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               )                    �?��=��?�            Pt@               (                   �a@�q�q�?             >@              !                    �?�eP*L��?             6@                                   �P@�q�q�?             (@                                  �?z�G�z�?             $@                                  �a@      �?             @        ������������������������       �                     �?                                  �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        "       %                 ����?z�G�z�?             $@        #       $                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        &       '                   �U@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        *       e                    �?�
 �^�?�            pr@       +       b                   h@|0M�Y4�?�            �p@       ,       a       	             �?��ckݭ�?�            �p@       -       J                    �?���c���?d            �c@        .       E                 ����?���*�?)             N@       /       4                    T@��Sݭg�?            �C@        0       3                    �?�q�q�?             @       1       2                    пz�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        5       D                    �?"pc�
�?            �@@       6       ?                   �q@     ��?             @@       7       8                    �?�>����?             ;@        ������������������������       �                      @        9       >                   `i@�KM�]�?             3@        :       ;                 �����      �?             @        ������������������������       �                     �?        <       =                   @`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             .@        @       C                    �?���Q��?             @       A       B                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        F       I       
             �?���N8�?             5@        G       H                    �N@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        K       ^                   �b@8��8���?;             X@       L       M                   �b@��S�ۿ?7            �V@       ������������������������       �                     �I@        N       [                    �?8�Z$���?            �C@       O       Z                    p@<���D�?            �@@       P       Q                    �?"pc�
�?             6@        ������������������������       �                     @        R       W                   �m@���y4F�?             3@       S       V                   �_@��S�ۿ?	             .@       T       U                    �I@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        X       Y                    _@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        \       ]                   �O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        _       `                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        G            @[@        c       d                    d@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        f       o                    @K@r�q��?             8@        g       h                    \@      �?              @        ������������������������       �                     �?        i       n                    �?؇���X�?             @        j       m                   �d@      �?             @       k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        p       w                   @b@     ��?             0@       q       r                    �?8�Z$���?             *@        ������������������������       �                     �?        s       v                   �Y@�8��8��?
             (@        t       u                 `ff�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        y       �                   �a@*
;&���?�             w@        z       �                    �?�x�E~�?6            @V@        {       �                    `Q@���}<S�?             7@       |       }                 ����?���7�?             6@       ������������������������       �        	             ,@        ~                           �M@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        &            �P@        �       �                    �?�n`���?�            pq@        �       �                    �?�������?"             N@       �       �                   �b@��k��?            �J@       �       �                    �B@�q�q�?             E@        ������������������������       �                     @        �       �                    �?�d�����?             C@       �       �       
             �?�����?             5@        ������������������������       �                     @        �       �                    @H@�t����?
             1@        ������������������������       �                     @        �       �                 ����?"pc�
�?             &@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?��.k���?	             1@       �       �                    �O@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @H@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                    �B@���U@��?�            `k@        �       �                    �?����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?0��_��?�            �j@        �       �       	             �?d�;lr�?)            �O@       �       �                   �b@^�!~X�?!            �J@       �       �                   `c@ >�֕�?            �A@       �       �                    �N@      �?             @@       ������������������������       �                     6@        �       �                   �`@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �l@�E��ӭ�?             2@        �       �                     O@r�q��?             @       �       �                    �?�q�q�?             @       �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?���Q��?             $@       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@8����?c            �b@       �       �                 ����?`���i��?9             V@        �       �                   �e@@9G��?            �H@       �       �                   �[@@��8��?             H@        �       �                    �?؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                    �M@Xny��?*            �N@        �       �                 ��� @�X����?             6@       �       �                    �?j���� �?             1@       �       �                    @M@�q�q�?
             (@       �       �                    �?      �?              @       �       �                    ^@      �?             @        ������������������������       �                      @        �       �                    �?      �?             @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ����?      �?             @       �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �C@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B�  ��� ���?���o���?�y��!�?.�u�y�?8��18�?28��1�?ffffff�?333333�?۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�c�1Ƹ?�s�9��?�$I�$I�?�m۶m��?              �?F]t�E�?]t�E�?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �<�@�0�?d���<�?UUUUUU�?UUUUUU�?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�������?      �?      �?              �?      �?              �?      �?      �?                      �?              �?{>�e���?�i
��?P��9��?~�3���?ZK���v�?1��:kI�?;�;��?�;�;�?""""""�?wwwwww�?�|˷|��?�i�i�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        /�袋.�?F]t�E�?      �?      �?�Kh/��?h/�����?      �?        �k(���?(�����?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?      �?      �?              �?      �?                      �?              �?��y��y�?�a�a�?�q�q�?�q�q�?      �?                      �?      �?        �������?�������?�������?�?      �?        ;�;��?;�;��?|���?|���?/�袋.�?F]t�E�?      �?        6��P^C�?(������?�������?�?�������?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?                      �?      �?              �?              �?      �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        8��Moz�?���,d!�?p�\��?����G�?d!Y�B�?ӛ���7�?F]t�E�?�.�袋�?              �?      �?      �?              �?      �?              �?                      �?�c�1��?�9�s��?�������?�������?oe�Cj��?"5�x+��?UUUUUU�?UUUUUU�?              �?Cy�5��?y�5���?=��<���?�a�a�?      �?        <<<<<<�?�?      �?        /�袋.�?F]t�E�?      �?      �?      �?                      �?      �?        �������?�?�������?�������?      �?                      �?              �?F]t�E�?]t�E�?      �?                      �?              �?��QNG9�?��5�X�?�m۶m��?�$I�$I�?      �?                      �?�V�9�&�?"5�x+��?�eY�eY�?��i��i�?�	�[���?�}�	��?�A�A�?��+��+�?      �?      �?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        r�q��?�q�q�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�y���?`��c.�?F]t�E�?F]t�E�?9/���?������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?      �?                      �?�}�K�`�?C��6�S�?]t�E]�?�E]t��?ZZZZZZ�?�������?�������?�������?      �?      �?      �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?      �?      �?      �?      �?              �?      �?              �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJOy�qhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�+         X                    �?p�Vv���?�           ��@                                  I@����l�?�            `w@                                   �?Dc}h��?#             L@                                 �[@П[;U��?             =@        ������������������������       �                     @               	                 433�?\X��t�?             7@                                   @D@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        
                           �?"pc�
�?	             &@                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                   W@PN��T'�?             ;@        ������������������������       �                     �?                      
             �?ȵHPS!�?             :@                                 0`@�LQ�1	�?             7@                                 @b@�}�+r��?             3@       ������������������������       �        
             0@                                   ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               7                    �?�Y���?�            �s@                                   �L@��SПW�?�            �j@                                 �f@����?l            �e@       ������������������������       �        k            `e@        ������������������������       �                     �?        !       "                   ``@�T|n�q�?            �E@        ������������������������       �        
             0@        #       6                 033@������?             ;@       $       %                    �?r�q��?             8@        ������������������������       �                     &@        &       5                    �?�	j*D�?
             *@       '       0                    �?      �?	             (@       (       /                    �?      �?              @       )       *                    �?r�q��?             @        ������������������������       �                     �?        +       .                    �?z�G�z�?             @        ,       -                   pa@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        1       2                     O@      �?             @        ������������������������       �                     �?        3       4                 hff�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        8       I                    �?�/���?C            �Y@       9       B                    l@�<ݚ�?'             K@        :       ;                   �a@�û��|�?             7@        ������������������������       �                     $@        <       A                    _@�	j*D�?
             *@       =       >                    �?      �?              @        ������������������������       �                     @        ?       @                    ]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        C       D                    �M@��a�n`�?             ?@       ������������������������       �                     :@        E       F                    �?���Q��?             @        ������������������������       �                      @        G       H                    `P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       M                    �? \� ���?            �H@        K       L                    �R@ףp=
�?             4@       ������������������������       �                     2@        ������������������������       �                      @        N       W                 ����?J�8���?             =@       O       P                    �D@      �?	             4@        ������������������������       �                     @        Q       R                   @`@      �?             0@        ������������������������       �                     @        S       T                    �?�C��2(�?             &@        ������������������������       �                      @        U       V                     M@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        Y       �                   0f@<�Z��?�            �v@       Z       �                   p`@\�c;��?�            Pv@        [       �                    �?֞R!R��?g             f@       \       e                    �?�ˡ�5��?T            �a@        ]       ^                   `X@�X����?             6@        ������������������������       �                      @        _       `                    �?      �?             4@        ������������������������       �                      @        a       d                 033�?�q�q�?             (@       b       c                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        f       �                    �?��(\���?H             ^@       g       h                   �h@�ܸb���?3             W@        ������������������������       �                     ?@        i       t                    �?f>�cQ�?#            �N@        j       s                    `@�q�q�?             2@       k       p                    �?z�G�z�?	             .@       l       o       	             �?8�Z$���?             *@       m       n                   �l@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        q       r                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        u       z                    �?Du9iH��?            �E@        v       y                   �m@�X�<ݺ?             2@        w       x                    �H@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        {       �                   �\@HP�s��?             9@        |       }                    �?����X�?             @        ������������������������       �                     �?        ~                          0i@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     <@        �       �                    �?����X�?            �A@        ������������������������       �                     @        �       �                    @J@J�8���?             =@        �       �                   a@"pc�
�?             &@       ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?X�<ݚ�?
             2@       �       �                    @���!pc�?             &@       �       �                   �i@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �       	             �?P���Q�?q            �f@       �       �                   `f@h�|�6�?i            @e@       �       �                    �?F|/ߨ�?d            @d@       �       �                   a@ ��ʻ��?U             a@       ������������������������       �        D             ]@        �       �                   Pa@ףp=
�?             4@        ������������������������       �                     �?        �       �                   �b@�}�+r��?             3@       ������������������������       �        	             "@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                   0p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     Q@$�q-�?             :@       �       �                    �?`2U0*��?             9@        �       �                   pc@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     �?        �       �                    �?      �?              @        �       �                    a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�
  w
��,@�?�z�����?����=��?n�ʄm�?۶m۶m�?�$I�$I�?��=���?�{a���?              �?!Y�B�?��Moz��?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?              �?h/�����?&���^B�?      �?        �؉�؉�?��N��N�?Y�B��?��Moz��?(�����?�5��P�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?                      �?'oe�C�?e�Cj���?���o.��?��0�?�}A_��?�}A_�w?      �?                      �?���)k��?6eMYS��?      �?        B{	�%��?{	�%���?�������?UUUUUU�?      �?        vb'vb'�?;�;��?      �?      �?      �?      �?�������?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��`����?�">�Tr�?9��8���?�q�q�?8��Moz�?��,d!�?      �?        ;�;��?vb'vb'�?      �?      �?      �?        �������?�������?              �?      �?                      �?�s�9��?�c�1Ƹ?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        և���X�?
^N��)�?�������?�������?              �?      �?        |a���?�rO#,��?      �?      �?              �?      �?      �?              �?]t�E�?F]t�E�?      �?        �q�q�?�q�q�?      �?                      �?              �?�[�[�?�>�>��?���վ?�I%�I%�?�L;k��?�,1>e��?H���@��?�RO�o��?�E]t��?]t�E]�?              �?      �?      �?      �?        �������?�������?      �?      �?      �?                      �?              �?333333�?�������?��,d!�?Nozӛ��?              �?�u�y���?��!XG�?UUUUUU�?UUUUUU�?�������?�������?;�;��?;�;��?      �?      �?      �?                      �?              �?      �?      �?              �?      �?              �?        w�qGܱ?qG�w��?�q�q�?��8��8�?�$I�$I�?۶m۶m�?      �?                      �?              �?{�G�z�?q=
ףp�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�$I�$I�?�m۶m��?              �?|a���?�rO#,��?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?r�q��?F]t�E�?t�E]t�?      �?      �?              �?      �?              �?                      �?�������?ffffff�?�?�������?�����H�?�Hx�5�?�?�������?              �?�������?�������?      �?        (�����?�5��P�?              �?�������?�������?              �?UUUUUU�?�������?              �?      �?        ;�;��?�؉�؉�?{�G�z�?���Q��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?              �?�������?�������?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��ghG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK݅�h��B@7         �                    �?.��X~��?�           ��@                                 �x@�Z���Z�?           �y@                                  �?���,_��?            �y@                                pff�?N1���?&            �N@                                 �r@`�(c�?            �H@                                 �b@�X����?             F@                                  �?���y4F�?             C@                               ����?r�q��?             B@       	       
                    [@      �?             8@        ������������������������       �                     @                                  �a@ףp=
�?             4@                                  `k@����X�?             @        ������������������������       �                     @                                  �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?      �?	             (@        ������������������������       �                     @        ������������������������       �                     "@                                  �U@@~�5��?�            �u@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               ~                    �R@�ʈD��?�            �u@              K                    �?lR���?�            pu@               F                   @e@��zi��?9            �V@               5       
             �?,�"���?6            @U@        !       *                   d@��P���?            �D@       "       )                 hff�?��a�n`�?             ?@        #       &                   �`@�θ�?             *@        $       %                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        '       (                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             2@        +       4                   �`@���Q��?             $@       ,       3                 033@      �?              @       -       .                   Pl@؇���X�?             @        ������������������������       �                     @        /       0                    �?      �?             @        ������������������������       �                      @        1       2                     J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        6       =                   �l@�C��2(�?             F@       7       8                    �?(;L]n�?             >@       ������������������������       �                     3@        9       <                    @K@�C��2(�?             &@        :       ;                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        >       ?                   �`@d}h���?
             ,@        ������������������������       �                     "@        @       A                     L@���Q��?             @        ������������������������       �                     �?        B       E                    �?      �?             @        C       D                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        G       H                    �?      �?             @        ������������������������       �                      @        I       J                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        L       }                   �a@(�s���?�            �o@       M       p                   pb@\� ���?w            �h@       N       [                    @L@ >�֕�?h            �e@       O       P                    @J@��:�-�?;            @Y@       ������������������������       �                     �I@        Q       X                    �?`2U0*��?             I@       R       W                   �[@��Y��]�?            �D@        S       T                   `[@��S�ۿ?	             .@       ������������������������       �                     (@        U       V                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        Y       Z                    �J@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        \       o                   �`@������?-            �R@       ]       n                   `@�㙢�c�?             G@       ^       k                   `_@r֛w���?             ?@       _       d                   �d@�J�4�?             9@       `       a                    �?      �?             0@       ������������������������       �                     ,@        b       c                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       j                    �?�q�q�?             "@       f       g                    _@և���X�?             @        ������������������������       �                     @        h       i                   �[@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             .@        ������������������������       �                     <@        q       r                     E@���N8�?             5@        ������������������������       �                      @        s       |                    �?�n_Y�K�?             *@       t       {                    �?���!pc�?	             &@       u       z                    �?և���X�?             @       v       w                   pd@���Q��?             @        ������������������������       �                      @        x       y                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        '             L@        ������������������������       �                     �?        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?T��ٟK�?�            �s@       �       �                    �?n�3���?�             s@       �       �                    �?LK�?.�?�            �p@       �       �                   @g@p=
ףp�?�             n@       �       �                    X@`.��A��?�            �m@        �       �                   �[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                     R@(.��H�?�            `m@       �       �                    @��xJ_�?�             m@       �       �       	             �?�NI���?�             m@       �       �                    P@     ��?I             `@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�-���e�?G            �_@        ������������������������       �                    �B@        �       �                    �?xP�Fֺ�?2            @V@       �       �                   �s@���?*            �R@       �       �                   �b@0�й���?)            @R@       ������������������������       �                    �C@        �       �                 ����?�������?             A@       �       �       
             �?�z�G��?             >@        �       �                   l@���|���?             &@       �       �                     E@      �?              @        ������������������������       �                     @        �       �                   `]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�KM�]�?	             3@       �       �                   0n@�t����?             1@       ������������������������       �                     ,@        �       �                   @[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        �       �                   0p@��9J���?C             Z@       ������������������������       �        *            @P@        �       �                   �?$�q-�?            �C@       ������������������������       �                     A@        �       �                    q@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `ff�?�g�y��?             ?@       �       �       
             �?�X����?             6@       �       �                    �?p�ݯ��?             3@       �       �                   `b@�q�q�?             (@       �       �                    @M@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    V@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�'�=z��?            �@@        ������������������������       �                     "@        �       �                    �?�q�q�?             8@        ������������������������       �                      @        �       �                   ``@�GN�z�?             6@        ������������������������       �                      @        �       �                   �c@X�Cc�?
             ,@       �       �                    �?�eP*L��?             &@       �       �                   �a@���Q��?             $@        �       �                    �?      �?             @       �       �                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �d@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@�q�q�?	             .@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �                   h@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��� ���?���o���?�G�5�?`�¼r�?�?�������?�:ڼO�?�}�K�`�?������?4և����?�E]t��?]t�E]�?6��P^C�?(������?�������?UUUUUU�?      �?      �?              �?�������?�������?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?      �?              �?                      �?              �?              �?      �?      �?      �?                      �?$�qe�?[̱]S��?UUUUUU�?UUUUUU�?              �?      �?        �}A_з?A_���?�|�&#�?k&{��?h�h��?��_��_�?�������?�?�����?������?�c�1Ƹ?�s�9��?�؉�؉�?ى�؉��?�������?333333�?              �?      �?              �?      �?      �?                      �?              �?333333�?�������?      �?      �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?      �?              �?      �?                      �?              �?F]t�E�?]t�E�?�?�������?              �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?۶m۶m�?I�$I�$�?              �?333333�?�������?              �?      �?      �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?��y��y�?�a�a�?������?c}h���?�A�A�?��+��+�?��be�F�?0��<�]�?              �?{�G�z�?���Q��?������?8��18�?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?�q�q�?      �?                      �?к����?��g�`��?d!Y�B�?�7��Mo�?�B!��?���{��?{�G�z�?�z�G��?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?��y��y�?�a�a�?              �?ى�؉��?;�;��?t�E]t�?F]t�E�?۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?                      �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?e�}��?�k���?�5��P�?�k(����?-0c����?K?s�y�?333333�?ffffff�?xp�zR�?@|4!/l�?      �?      �?              �?      �?        ç����?��jZǛ�?�k�u��?����S��?��FX��?���=��?      �?      �?      �?      �?      �?                      �?M�4M�4�?�eY�eY�?      �?        �.p��?�я~���?O贁N�?ƒ_,���?����?����Ǐ�?      �?        �������?�������?ffffff�?333333�?F]t�E�?]t�E]�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �k(���?(�����?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?      �?        ;�;��?�؉�؉�?      �?        �؉�؉�?;�;��?      �?        �������?333333�?              �?      �?                      �?              �?              �?��{���?�B!��?�E]t��?]t�E]�?^Cy�5�?Cy�5��?�������?�������?9��8���?�q�q�?      �?                      �?              �?�m۶m��?�$I�$I�?              �?      �?              �?                      �?|���?|��|�?      �?        �������?�������?      �?        ]t�E�?�袋.��?              �?�m۶m��?%I�$I��?]t�E�?t�E]t�?�������?333333�?      �?      �?      �?      �?              �?      �?              �?        UUUUUU�?�������?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?        �q�q�?r�q��?      �?        UUUUUU�?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJiƋ.hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�7         �                    �?�ܲ�}��?�           ��@              i                    �?j:?���?           �y@              T                   �b@,���i�?�            �t@                                  �?\E�w���?�            `r@                                   x@�q�q�?             8@                                   O@�㙢�c�?             7@       ������������������������       �                     (@                                   �?���|���?             &@       	       
                 `ff @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?               S                    �?�:�^���?�            �p@              2                   `_@H�g�}N�?v            �f@                                 `[@�o�s(��?J            �[@                                   �?�?�|�?            �B@                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ?@               #                    �?�F��O�?0            @R@               "                 pff�?z�G�z�?             .@              !                 ����?      �?              @                                 �]@����X�?             @        ������������������������       �                     @                       
             �?�q�q�?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        $       %                   `l@�8���?$             M@       ������������������������       �                     =@        &       -                    �?ܷ��?��?             =@        '       (                    @N@ףp=
�?             $@        ������������������������       �                     @        )       ,                    �O@z�G�z�?             @       *       +                   Pr@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        .       /                     K@�KM�]�?
             3@       ������������������������       �                     .@        0       1                    ]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        3       J       	             �?<ݚ�?,             R@       4       I                   �m@     ��?&             P@       5       H                   �m@�4F����?            �D@       6       ?                    �?�d�����?             C@        7       8                   �`@և���X�?             ,@        ������������������������       �                     @        9       >                   �h@z�G�z�?             $@        :       =                   @e@���Q��?             @       ;       <                   �g@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        @       C                   �_@r�q��?             8@        A       B                   �j@      �?             @        ������������������������       �                      @        ������������������������       �                      @        D       G                   P`@ףp=
�?             4@        E       F                   @_@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     7@        K       L                    �?      �?              @        ������������������������       �                      @        M       R                    �H@�q�q�?             @       N       Q                    �?�q�q�?             @       O       P                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        2             V@        U       Z                 ����?�!���?             A@        V       W                     G@      �?              @        ������������������������       �                     @        X       Y                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        [       f                    �?�n_Y�K�?             :@       \       e                    @N@�\��N��?             3@       ]       d                    @     ��?             0@       ^       a                    �?���Q��?
             .@       _       `                   ``@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        b       c                   @`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        g       h                    @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        j              
             �?>���Rp�?2            �U@       k       ~                    �?�Y����?(            �P@        l       y                    �?���@M^�?             ?@       m       x                 833@
j*D>�?             :@       n       u       	             �?b�2�tk�?             2@       o       r                    �?���Q��?             $@        p       q                   �t@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        s       t                   p@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        v       w                    @L@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        z       {                   P`@z�G�z�?             @        ������������������������       �                      @        |       }                   c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     B@        �       �                    �?�G�z��?
             4@        ������������������������       �                     @        �       �                 ����?8�Z$���?             *@       �       �                   �b@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   `_@h
WY�v�?�            �s@        �       �                    �I@"Ae���?            �G@        �       �                    �E@�����?             5@        �       �                   �]@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             1@        �       �                    ^@��
ц��?             :@       �       �                    �?������?
             .@        ������������������������       �                     @        �       �                   @V@      �?              @        ������������������������       �                     �?        �       �                    �?և���X�?             @        �       �                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @33�?      �?             @       �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `c@�C��2(�?             &@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�G�V�e�?�             q@       �       �                 ���@�mm�y��?�            @o@       �       �                    @M@��a_�U�?�            `n@       �       �                   @g@�qW$�a�?z            `i@       �       �                   �O@�G� �?y            @i@        ������������������������       �                     �?        �       �                    �?0�,���?x             i@       �       �                 ����?@3�qH�?a             d@       �       �                    �?���б�?P            �`@        ������������������������       �                     =@        �       �                    �?@䯦s#�?=            �Z@       �       �       
             �?�����?:            @Y@       ������������������������       �        &            @Q@        �       �                   �c@      �?             @@        �       �                   �b@      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        ������������������������       �        
             0@        ������������������������       �                     @        ������������������������       �                     :@        �       �                    �?      �?             D@       �       �                   xq@r�q��?             >@       �       �                    �?���}<S�?             7@       �       �                    @D@�}�+r��?             3@        �       �                   �e@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        �       �                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Xr@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    ]@�z�G��?             D@        �       �                   �a@�q�q�?             @        ������������������������       �                     @        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@������?             A@       ������������������������       �                     6@        �       �       	             �?�q�q�?             (@       �       �                    r@���!pc�?             &@       �       �                   �i@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   hq@8�A�0��?             6@       �       �                   �j@z�G�z�?
             .@        �       �                    a@      �?             @       �       �                   @`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ����u��?/�E��?e��N���?'�B��K�?8��18�?�����?P&�to@�?6;j���?�������?UUUUUU�?d!Y�B�?�7��Mo�?              �?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?              �?      �?              �?      �?      �?                      �?      �?        l�l��?}�'}�'�?���?|��{���?J��yJ�?�k߰��?к����?*�Y7�"�?UUUUUU�?�������?      �?                      �?              �?�P�B�
�?�իW�^�?�������?�������?      �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?                      �?a���{�?j��FX�?              �?a���{�?��=���?�������?�������?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?(�����?�k(���?              �?      �?      �?      �?                      �?��8��8�?�q�q�?      �?     ��?KԮD�J�?ە�]���?y�5���?Cy�5��?۶m۶m�?�$I�$I�?      �?        �������?�������?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?�������?      �?      �?      �?                      �?�������?�������?�q�q�?9��8���?              �?      �?                      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?�������?�������?      �?      �?              �?      �?      �?              �?      �?        ى�؉��?;�;��?�5��P�?y�5���?      �?      �?333333�?�������?]t�E]�?F]t�E�?      �?                      �?      �?      �?              �?      �?                      �?              �?�$I�$I�?۶m۶m�?              �?      �?        GX�i���?�i��F�?���@���?��¯�D�?�c�1��?�s�9��?;�;��?b'vb'v�?�8��8��?9��8���?333333�?�������?�������?333333�?              �?      �?        �������?�������?      �?                      �?      �?      �?      �?                      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?        ;�;��?;�;��?�$I�$I�?�m۶m��?              �?      �?                      �?��f����?�e�}��?�w6�;�?W�+���?=��<���?�a�a�?      �?      �?      �?                      �?      �?        �؉�؉�?�;�;�?wwwwww�?�?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?                      �?              �?F]t�E�?]t�E�?�������?�������?      �?                      �?              �?�������?�������?%��C��?���S㥻?�����]�?;����?���)��?��%f-�?�tj��?�~�X��?              �?Ez�rv�?g��1��?��6��?r���py?5�m�Q��?t��:W~?      �?        R����?�x+�R�?�tj��?��be�F�?      �?              �?      �?      �?      �?      �?                      �?      �?              �?              �?              �?      �?�������?UUUUUU�?ӛ���7�?d!Y�B�?�5��P�?(�����?�������?�������?      �?                      �?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?                      �?ffffff�?333333�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?xxxxxx�?�?      �?        UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?333333�?�������?              �?      �?                      �?      �?                      �?颋.���?/�袋.�?�������?�������?      �?      �?      �?      �?              �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ*�/shG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK녔h��B�:         f                 033�?�ܲ�}��?�           ��@              7                    �?rLB0J-�?�            �w@                                 �c@0������?�            @n@                                ����?
j*D>�?             :@                                  @J@r�q��?             2@                                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        	                           �?$�q-�?             *@        
                           ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @               "                    �?d/
k�?�             k@              !       	             �?0m��5!�?p            �f@                                  @t@�IєX�?,             Q@                                  @G@�g�y��?)             O@        ������������������������       �                     ;@                                   �G@ >�֕�?            �A@                                  �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �i@Pa�	�?            �@@                                  @i@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@                                 ����?�q�q�?             @                                  �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        D            @\@        #       4                    �?��
P��?            �A@       $       /                 ����?l��[B��?             =@       %       .                    �?�����?             3@       &       -                   �c@      �?             (@       '       ,                    �?�q�q�?             "@       (       +                    �?؇���X�?             @       )       *                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        0       1                    @M@ףp=
�?             $@       ������������������������       �                      @        2       3                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       6                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        8       C                    �?N�Q�z��?_             a@       9       :                   �g@ДX��?0             Q@        ������������������������       �                     @@        ;       <                    �I@tk~X��?             B@        ������������������������       �                     0@        =       B                    �?��Q��?             4@       >       ?                 ����?���|���?	             &@        ������������������������       �                     @        @       A                    b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        D       I                    @D@bKv���?/            @Q@        E       F                   @d@�C��2(�?             &@       ������������������������       �                     @        G       H                    a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        J       K                   @[@�c�Α�?*             M@        ������������������������       �                     @        L       Q                   @E@l��
I��?(             K@        M       N                   @_@����X�?             @        ������������������������       �                     @        O       P                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        R       W                   �c@��|�5��?#            �G@       S       V                    `P@      �?             @@       T       U                    �?��S�ۿ?             >@       ������������������������       �                     <@        ������������������������       �                      @        ������������������������       �                      @        X       ]                    �?��S���?             .@        Y       \                    �?z�G�z�?             @       Z       [                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ^       e                 @33�?���Q��?	             $@       _       `                   �i@X�<ݚ�?             "@        ������������������������       �                     @        a       d                   �d@z�G�z�?             @        b       c                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        g       �                    �?�j����?�            0v@       h       �                   �c@�m�6�?�             s@       i       �                    �?�&�F��?�            �p@        j       q                    �?      �?'             J@        k       p       	             �?��2(&�?             6@       l       m                    �Q@r�q��?             2@       ������������������������       �                     ,@        n       o                 hff@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        r       �                   �p@�q�q�?             >@       s       v                    �?      �?             8@        t       u                   @\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        w       x                    @F@���N8�?             5@        ������������������������       �                     @        y       z                   Pm@�����H�?             2@       ������������������������       �                     $@        {       �                    �?      �?              @       |       }                    �?؇���X�?             @       ������������������������       �                     @        ~                          `@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@�q�q�?             @        ������������������������       �                     @        �       �       	             �?�q�q�?             @       �       �                   `^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��<nd�?�            @k@        �       �                    S@� ��1�?            �D@        ������������������������       �                     �?        �       �                    �?z�G�z�?             D@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �R@�t����?             A@       �       �                    �?      �?             @@        ������������������������       �        
             ,@        �       �                   �W@�����H�?
             2@        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                      @        �       �                   Pr@�O2�J�?o             f@       �       �                   0j@X�.�d�?[            �a@        �       �                    b@ ,��-�?'            �M@       �       �                   �i@ ��WV�?#             J@       �       �                   ``@@�E�x�?!            �H@       �       �                    �?���N8�?             5@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     <@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �b@����X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��'�`�?4            �T@       �       �                   8p@�k~X��?-             R@       ������������������������       �                     H@        �       �                    �? �q�q�?             8@       ������������������������       �                     4@        �       �                   `\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                 ����?؇���X�?            �A@        �       �                    �?     ��?             0@       �       �                    �?r�q��?             (@       �       �                    @I@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    [@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        �       �       
             �?      �?             B@       �       �       	             �?��H�}�?             9@       �       �                   �r@r�q��?	             (@       ������������������������       �                     $@        ������������������������       �                      @        �       �                   �d@��
ц��?             *@       �       �                   d@���|���?             &@       �       �                    @H@�q�q�?             @       �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                     J@"pc�
�?             &@        ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                    U@�`���?             �H@        �       �                    �?�t����?	             1@        ������������������������       �                     @        �       �                 `ff�?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �                    r@     ��?             @@       �       �                    �?�+e�X�?             9@       �       �                 ���@�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        �       �                    �?      �?              @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?և���X�?             @       �       �                   �\@      �?             @        ������������������������       �                      @        �       �                    �H@      �?             @        ������������������������       �                      @        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �t�b�`     h�h)h,K ��h.��R�(KK�KK��hi�B�  ����u��?/�E��?ި2�ć�?E���v��?�V���?������?;�;��?b'vb'v�?UUUUUU�?�������?�������?333333�?              �?      �?        ;�;��?�؉�؉�?      �?      �?      �?                      �?              �?      �?        �Kh/���?/�����?kdu�J�?�rS�<��?�?�?��{���?�B!��?      �?        ��+��+�?�A�A�?      �?      �?              �?      �?        |���?|���?۶m۶m�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        _�_��?PuPu�?���=��?GX�i���?^Cy�5�?Q^Cy��?      �?      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?              �?                      �?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        )�[�?r��8R�?ZZZZZZ�?�������?              �?9��8���?r�q��?              �?ffffff�?�������?]t�E]�?F]t�E�?              �?      �?      �?      �?                      �?              �??���(��?��v`��?F]t�E�?]t�E�?              �?UUUUUU�?�������?      �?                      �?5�rO#,�?�{a���?      �?        Lh/����?h/�����?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?        br1���?x6�;��?      �?      �?�������?�?      �?                      �?              �?�?�������?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?333333�?�q�q�?r�q��?              �?�������?�������?      �?      �?      �?                      �?      �?                      �?z}]5R�?�`��rk�?�)�)�?�5��5��?Hֹ�d�?7Ũ�oS�?      �?      �?t�E]t�?��.���?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        ��y��y�?�a�a�?      �?        �q�q�?�q�q�?              �?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?4R1�:#�?����[�?������?������?      �?        ffffff�?ffffff�?      �?      �?              �?      �?        �?<<<<<<�?      �?      �?              �?�q�q�?�q�q�?      �?                      �?      �?        k��2�?�v�,1�?�@�6�?�ۥ����?'u_[�?[4���?;�;��?O��N���?9/���?և���X�?�a�a�?��y��y�?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?��k���?1P�M��?�q�q�?�8��8��?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?�������?�������?�������?      �?                      �?              �?      �?      �?              �?      �?                      �?      �?      �?
ףp=
�?{�G�z�?UUUUUU�?�������?              �?      �?        �;�;�?�؉�؉�?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?/�袋.�?F]t�E�?      �?        333333�?�������?              �?      �?        և���X�?����S�?�?<<<<<<�?              �?F]t�E�?/�袋.�?              �?      �?              �?      �?R���Q�?���Q��?�?�?      �?                      �?      �?      �?      �?      �?      �?              �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��\hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         �                    �?8}�ý�?�           ��@              E                    �?��Sz�?	           �z@                                  �?������?�            �q@                      	             �?      �?
             2@                                  �?X�Cc�?             ,@                                  �?�eP*L��?             &@                                  �?�q�q�?             "@        ������������������������       �                      @        	       
                   `\@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               D                 ���@8Ӈ���?�            `p@              9                    �?�:�]��?�            �o@              ,                    �?�2�~w�?�            �k@                                  �?蹱f
@�?i            �e@                               pff�?@	tbA@�?Q            @a@                     
             �?�Ru߬Α?E            �\@       ������������������������       �        /            �S@                                  @t@������?             B@       ������������������������       �                    �A@        ������������������������       �                     �?                                   �? �q�q�?             8@       ������������������������       �                     1@                                   a@؇���X�?             @                                  �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                !                    U@z�G�z�?            �A@        ������������������������       �                     @        "       +                   pf@      �?             @@       #       (                   �o@��S�ۿ?             >@       $       %                    b@ �q�q�?             8@       ������������������������       �                     5@        &       '                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        )       *                    �K@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        -       6                   �?dP-���?            �G@       .       /                    迀��7�?             F@        ������������������������       �                     �?        0       5                    T@ qP��B�?            �E@        1       2                    �?؇���X�?             @        ������������������������       �                     @        3       4                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     B@        7       8                   @c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        :       ;                    �?z�G�z�?            �A@        ������������������������       �                     .@        <       ?                    �?��Q��?             4@        =       >                   �b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        @       A                   �b@���Q��?             $@        ������������������������       �                      @        B       C                   �f@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        F       Y                    �?����*�?`             b@        G       H                   �Q@�c�Α�?             =@        ������������������������       �                     @        I       R                    �?���B���?             :@       J       K                 ����?�t����?             1@        ������������������������       �                     @        L       M                   `X@z�G�z�?	             $@        ������������������������       �                     �?        N       Q                    @J@�����H�?             "@        O       P                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        S       X                 ����?�q�q�?             "@       T       U                 ����?؇���X�?             @        ������������������������       �                     @        V       W                    b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        Z       u                    �?Riv����?I             ]@        [       r                    �?�q����?!            �J@       \       m                   0a@�ʻ����?             A@       ]       f                   �_@�û��|�?             7@       ^       e                   pf@��S���?	             .@       _       `                    ]@�q�q�?             (@        ������������������������       �                     @        a       d                    @M@և���X�?             @       b       c                 ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        g       l                    �?      �?              @       h       i                   �`@r�q��?             @        ������������������������       �                     @        j       k       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        n       o                    �?�C��2(�?             &@       ������������������������       �                      @        p       q                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        s       t                     Q@�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        v       w                   �_@�i�y�?(            �O@        ������������������������       �                     A@        x       �                    �? 	��p�?             =@       y       |                    �?�t����?             1@        z       {                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        }       ~                   a@�C��2(�?             &@       ������������������������       �                     @               �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             (@        �       �                    V@�v�G���?�            Ps@        ������������������������       �                     @        �       �                    �?R��Xp�?�             s@        �       �                   �`@��.k���?             A@        �       �                    �?�q�q�?             2@        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @J@������?	             .@        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             0@        ������������������������       �                     @        �       �                    �L@X�<ݚ�?             "@       �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�Aʑ���?�            �p@       �       �                   Pb@ ���]��?�            �p@       �       �                    �?`�q��־?�             m@       �       �                   �e@h�����?p            `f@       �       �                    �?������?o            @f@       �       �                    �L@��F��?d            `c@       �       �                   `_@�ʈD��?8            �U@       �       �                   �[@��GEI_�?)            �N@        �       �                   �Z@؇���X�?             <@       �       �                    @L@�C��2(�?             6@       ������������������������       �        
             1@        �       �                   �a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �@@        �       �                   �_@�J�4�?             9@        �       �                 033@և���X�?             @       �       �                 ����?���Q��?             @        ������������������������       �                     �?        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �m@�X�<ݺ?             2@        ������������������������       �                     "@        �       �                   �^@�����H�?             "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        ,            @Q@        �       �                    �?��+7��?             7@       �       �                 `ff�?ҳ�wY;�?             1@       �       �                   0a@8�Z$���?             *@        ������������������������       �                     @        �       �                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     K@        �       �                    �?�4�����?             ?@        �       �                   �b@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �Z@��<b���?             7@        ������������������������       �                     @        �       �                   �d@ףp=
�?             4@       ������������������������       �        	             1@        �       �                     K@�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  a[ӿc�?PR Np�?O���N�?b���.b�?,��+���?PuPu�?      �?      �?�m۶m��?%I�$I��?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?                      �?      �?        �*NHɳ�?����a�?}}}}}}�?�?־a��?A��)A�?Z/`��U�?\
�IƢ�?�%~F��?ہ�v`��?���#��?p�}��?      �?        �q�q�?�q�q�?      �?                      �?�������?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?      �?      �?�������?�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?                      �?              �?�����F�?W�+�ɵ?�.�袋�?F]t�E�?              �?��}A�?�}A_З?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?        �������?ffffff�?�������?�������?      �?                      �?�������?333333�?      �?              �?      �?              �?      �?                      �?�k%�6�?'Jvm�d�?5�rO#,�?�{a���?              �?��؉���?ى�؉��?<<<<<<�?�?      �?        �������?�������?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?	�=����?>�����?�x+�R�?�Cj��V�?<<<<<<�?�������?8��Moz�?��,d!�?�������?�?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?      �?              �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?      �?        (�����?�5��P�?              �?      �?        AA�?�������?              �?�{a���?������?�?<<<<<<�?UUUUUU�?�������?              �?      �?        F]t�E�?]t�E�?              �?      �?      �?      �?                      �?              �?��O �?C���?      �?        �5��P^�?���k(�?�������?�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �?wwwwww�?      �?      �?      �?                      �?              �?      �?      �?      �?        r�q��?�q�q�?�������?UUUUUU�?      �?        �������?�������?              �?      �?                      �?Ũ�oS��?���u��?>���>�?���>��?r؃H{�?��6���?J���s�?wn�Q�?B�P�"�?ؽ�u�{�?mЦm�?Y���/Y�?�}A_з?A_���?;ڼOqɰ?�d����?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?              �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?{�G�z�?�z�G��?۶m۶m�?�$I�$I�?333333�?�������?              �?      �?      �?      �?                      �?              �?�q�q�?��8��8�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?              �?Y�B��?zӛ����?�������?�������?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?                      �?��RJ)��?���Zk��?      �?      �?              �?      �?        ��Moz��?��,d!�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKх�h��B@4         h                    �K@�/�$�y�?�           ��@              %                    �?ڬ`Z�s�?           Py@                                   �?*K�U��?�            `j@                                  I@Ћ����?g            �d@                                   �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                  h@`�V���?c            �c@       	       
       
             �?@f����?b            �c@       ������������������������       �        9            @V@                                  @[@�\=lf�?)            �P@                                   �?�q�q�?             @                                 �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        &             P@        ������������������������       �                     �?               $                    �?�[�IJ�?            �G@                                  �?X�<ݚ�?            �F@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                  �p@^H���+�?            �B@                                 �`@     ��?             @@                                  �?�ՙ/�?             5@        ������������������������       �                      @        ������������������������       �                     *@                                  b@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                !                    �H@z�G�z�?             @        ������������������������       �                      @        "       #                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        &       a                    �?��B���?�            @h@       '       H                    �I@�q�q�?e             b@       (       )                    @C@k�q��?=            @U@        ������������������������       �                     "@        *       9                    �?:W��S��?7             S@       +       2                   �m@��P���?            �D@       ,       -                 033@�C��2(�?             6@       ������������������������       �                     2@        .       1                    �?      �?             @       /       0                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        3       8                   �b@p�ݯ��?             3@       4       7                   @_@$�q-�?             *@        5       6                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             "@        ������������������������       �                     @        :       G                    d@؇���X�?            �A@       ;       <                    �?�GN�z�?             6@        ������������������������       �                     @        =       D                    �?�E��ӭ�?             2@       >       C                    �?���!pc�?             &@       ?       B                    @H@z�G�z�?             $@       @       A                     E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        E       F                 hff�?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             *@        I       N                    �?@�r-��?(            �M@        J       K                   �`@���Q��?             $@        ������������������������       �                     @        L       M                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        O       `                   pp@��<D�m�?             �H@       P       U                    @J@�L���?            �B@        Q       T                    b@z�G�z�?             @        R       S                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        V       Y                    �?      �?             @@        W       X                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        Z       _                   �[@`2U0*��?             9@        [       ^                    �?ףp=
�?             $@        \       ]                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �        	             (@        b       g                    �? "��u�?             I@       c       f                    �?ܷ��?��?             =@        d       e                   `\@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             4@        ������������������������       �                     5@        i       �                 pff�?�7����?�            �t@        j                           �?4ʟ����?O            �]@       k       |                   Pt@8^s]e�?)             M@       l       w                   �c@Ȩ�I��?'            �J@       m       p                    �?�3Ea�$�?"             G@        n       o                   �a@��
ц��?	             *@       ������������������������       �                     @        ������������������������       �                     @        q       r       	             �?�FVQ&�?            �@@       ������������������������       �                     0@        s       v                     M@�t����?             1@        t       u                    @L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             (@        x       {                   �]@����X�?             @        y       z                    Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        }       ~                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pb@�-ῃ�?&            �N@        ������������������������       �                     4@        �       �                 ����?D^��#��?            �D@       �       �                    �?��>4և�?             <@        �       �                    d@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���N8�?             5@       �       �                    �?�n_Y�K�?	             *@        ������������������������       �                     @        �       �                    �N@      �?              @       �       �                   Pp@և���X�?             @       �       �                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?8�Z$���?             *@        �       �                   �a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �R@�r�.kx�?�            @j@       �       �                   �`@�d2 Λ�?�            �i@        �       �                    `@�4���L�?8            �U@       �       �                    �P@(��+�?'            �N@       �       �                    �?�j��b�?%            �M@       �       �                    �?�S����?             C@       �       �                 `ff�?�����H�?             B@        �       �                   �^@�θ�?	             *@       �       �                    �L@r�q��?             (@        �       �                   �\@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    [@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                      @        �       �                    �?��H�}�?             9@        ������������������������       �                     @        �       �                   @X@���N8�?             5@        �       �                    �M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   r@      �?             0@       ������������������������       �                     &@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����˵�?M            �]@        �       �                   8t@�㙢�c�?             7@       �       �                    �?��2(&�?             6@       �       �                    �?      �?             0@        �       �                    j@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                     N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    a@ r���?;            �W@       ������������������������       �        -             Q@        �       �                    �?�>����?             ;@        ������������������������       �                     &@        �       �                    �?      �?	             0@       �       �                    d@�<ݚ�?             "@       �       �                    �?      �?              @       ������������������������       �                     @        �       �                    n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B  L�f���?Z�L��?+̉�?�g�����? � g���?��|c��?ԮD�J��?��+Q��?۶m۶m�?�$I�$I�?      �?                      �?�����?Kz���?�|˷|��?�A�Az?      �?        "=P9���?g��1��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?                      �?m�w6�;�?���
b�?�q�q�?r�q��?      �?      �?              �?      �?        �g�`�|�?L�Ϻ��?      �?      �?�a�a�?�<��<��?      �?                      �?F]t�E�?]t�E�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?��,O"��?(�i�n��?UUUUUU�?UUUUUU�?]]]]]]�?QQQQQQ�?              �?����k�?���k(�?�����?������?F]t�E�?]t�E�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?Cy�5��?^Cy�5�?;�;��?�؉�؉�?      �?      �?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?�袋.��?]t�E�?      �?        �q�q�?r�q��?F]t�E�?t�E]t�?�������?�������?      �?      �?      �?                      �?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?      �?        ��c+���?'u_�?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?և���X�?��S�r
�?L�Ϻ��?}���g�?�������?�������?      �?      �?      �?                      �?              �?      �?      �?�$I�$I�?۶m۶m�?              �?      �?        {�G�z�?���Q��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?���Q��?�G�z�?a���{�?��=���?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?G}g����?]AL� &�?�����?_̧^̧�?|a���?	�=����?+�R��?�	�[���?����7��?��,d!�?�؉�؉�?�;�;�?              �?      �?        >����?|���?      �?        <<<<<<�?�?333333�?�������?      �?                      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?                      �?�����?�).�u�?              �?,Q��+�?�]�ڕ��?I�$I�$�?۶m۶m�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��y��y�?�a�a�?ى�؉��?;�;��?              �?      �?      �?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?      �?                      �?;�;��?;�;��?333333�?�������?      �?                      �?      �?        �����?L��K���?�����ܼ?dddddd�?S֔5eM�?kʚ����?;ڼOq��?q�����?��/���?�N��?^Cy�5�?(������?�q�q�?�q�q�?�؉�؉�?ى�؉��?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        d!Y�B�?�Mozӛ�?      �?                      �?      �?                      �?      �?        
ףp=
�?{�G�z�?      �?        ��y��y�?�a�a�?�������?�������?      �?                      �?      �?      �?              �?�������?�������?      �?                      �?��/���?W'u_�?d!Y�B�?�7��Mo�?t�E]t�?��.���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �X�0Ҏ�?9�{n�S�?              �?h/�����?�Kh/��?              �?      �?      �?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJxS�ohG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKх�h��B@4         d                    �?�3u���?�           ��@                                  �?��G
L�?�            @w@               
                    �?�q�q��?             H@                                   �?���|���?             &@                                  @M@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?               	                    �G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                    K@������?            �B@        ������������������������       �                     �?                                   �?�8��8��?             B@                                  a@R���Q�?             4@                                  `^@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �        	             0@               U       	             �?����?�?�            @t@              <                 ����?�zӝ���?�            @i@              3                   �b@      �?a             c@              .                    �P@�O��/�?Y            `a@                                 �b@�U�=���?T            �`@       ������������������������       �        ,             R@                                  c@r�q��?(             N@        ������������������������       �                     @                                   �?���5��?'            �L@        ������������������������       �        
             0@               -                   0f@��r._�?            �D@              (                   �`@ �o_��?             9@                '                    �?և���X�?
             ,@       !       "                 ���ٿz�G�z�?             $@        ������������������������       �                     �?        #       &       
             �?�����H�?             "@        $       %                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        )       ,       
             �?�C��2(�?
             &@        *       +                   @j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@        /       2                    a@և���X�?             @       0       1                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        4       ;       
             �?�n_Y�K�?             *@       5       :                    �?X�<ݚ�?             "@       6       7                   �c@r�q��?             @        ������������������������       �                     @        8       9                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        =       >                    �?���Q��?%             I@        ������������������������       �                     @        ?       B                 `ff�?�X����?              F@        @       A       
             �?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        C       R                   q@�P�*�?             ?@       D       Q                   po@$��m��?             :@       E       P                   Pm@8�A�0��?             6@       F       I                    �?��Q��?             4@        G       H                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        J       O                    c@�t����?             1@       K       L                 033�?؇���X�?
             ,@       ������������������������       �                     $@        M       N                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        S       T                   �Z@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        V       _                    �? ;=֦��?L            �^@       W       X                    �?���͡?F            @\@        ������������������������       �                     >@        Y       Z                   �o@ Df@��?2            �T@       ������������������������       �                      K@        [       ^                   pg@ 	��p�?             =@       \       ]                   Xp@h�����?             <@        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                     �?        `       c                   @`@�����H�?             "@        a       b                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        e       �                   P`@��/�8�?�            �v@       f       �                 pff�?����?�            �i@       g       h                 ����?�$��y��?B            @X@        ������������������������       �                     G@        i       t                   �o@@�0�!��?#            �I@       j       m                    �?�C��2(�?            �@@        k       l                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        n       s                 033�? 	��p�?             =@        o       p                    �?�q�q�?             @        ������������������������       �                      @        q       r                   �[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        u       �                    �?�q�q�?             2@       v       y                   �Z@���Q��?
             .@        w       x                   �p@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        z       �       
             �?z�G�z�?             $@       {       |                    �?�����H�?             "@        ������������������������       �                     @        }       �                   �^@r�q��?             @        ~                           �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ]@����r�?A            �[@        �       �                   �[@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        =             Z@        �       �       	             �?���]�?a            `c@       �       �                    �?���4Z��?R            ``@       �       �                    �?��t���?6            �S@        �       �                 @33�?$��m��?             :@        ������������������������       �                     @        �       �                    �L@�G�z��?             4@       �       �                 ����?d}h���?
             ,@        �       �                    _@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    m@�C��2(�?             &@        ������������������������       �                     @        �       �                   @_@      �?             @        ������������������������       �                      @        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?0��_��?#            �J@       �       �                   �e@�ݜ�?            �C@       �       �                    �?�KM�]�?             C@        ������������������������       �                     "@        �       �                   ``@\-��p�?             =@        �       �                   @n@      �?	             (@        �       �                    �?      �?             @       �       �                    �F@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@�IєX�?	             1@       ������������������������       �                     (@        �       �                    @N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                    �?�n_Y�K�?             J@       �       �                    @J@v�X��?             F@        �       �                    �F@      �?             (@       �       �                    a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �Z@      �?             @@        ������������������������       �                     �?        �       �                   �c@��a�n`�?             ?@       �       �                   @p@`2U0*��?             9@       ������������������������       �        	             2@        �       �                   �p@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `t@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 lffֿ      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   d@�q�q�?             8@       �       �                 `ff�?X�<ݚ�?             2@       �       �                   �l@���|���?             &@        ������������������������       �                     @        �       �                    �?և���X�?             @       �       �                   �p@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    b@؇���X�?             @        �       �                 `ff�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B  k�w죻�?��	."�?X`�X�?�~�駟�?UUUUUU�?�������?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?      �?                      �?к����?��g�`��?      �?        UUUUUU�?UUUUUU�?333333�?333333�?t�E]t�?F]t�E�?      �?                      �?              �?              �?~X�<��?�n���?�(0��<�?�]?[��?      �?      �?*ۻ���?�&!��ȹ?�M6�d��?e�M6�d�?      �?        �������?UUUUUU�?              �?�}��?��Gp�?      �?        �ڕ�]��?ە�]���?
ףp=
�?�Q����?�$I�$I�?۶m۶m�?�������?�������?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        ;�;��?ى�؉��?�q�q�?r�q��?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?              �?        �������?333333�?      �?        ]t�E]�?�E]t��?;�;��?�؉�؉�?              �?      �?        �Zk����?�RJ)���?vb'vb'�?�N��N��?/�袋.�?颋.���?ffffff�?�������?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?              �?                      �?�������?�������?              �?      �?        �%C��6�?XG��).�?$��Co�?x�!���?      �?        c��7�:�?��k���?      �?        ������?�{a���?�m۶m��?�$I�$I�?              �?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?              �?        ӟ���?�8x��?ᖚ���?�V&O@t�?W?���?����?              �?�������?ZZZZZZ�?F]t�E�?]t�E�?      �?      �?      �?                      �?�{a���?������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?�������?�������?      �?                      �?�������?�������?�q�q�?�q�q�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?��)A��?�oX����?UUUUUU�?�������?              �?      �?                      �?�=���?�qa�?Ls�U��?ZF�ձ�?^-n����?�td�@T�?vb'vb'�?�N��N��?              �?�������?�������?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?]t�E�?              �?      �?      �?              �?      �?      �?      �?                      �?      �?        �V�9�&�?"5�x+��?�i�i�?\��[���?(�����?�k(���?              �?�{a���?a����?      �?      �?      �?      �?�������?333333�?              �?      �?              �?                      �?�?�?              �?�������?�������?      �?                      �?      �?                      �?ى�؉��?;�;��?颋.���?�.�袋�?      �?      �?      �?      �?      �?                      �?      �?              �?      �?      �?        �c�1Ƹ?�s�9��?{�G�z�?���Q��?              �?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �������?�������?�q�q�?r�q��?]t�E]�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?333333�?�������?              �?      �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQ ghG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�/         X                    �?�^�P��?�           ��@                                 �^@������?�            @x@                                   �?�!���?)             Q@                                  Z@�&!��?            �E@                                  �_@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @                                  `]@^H���+�?            �B@        	       
                    �?�C��2(�?             &@        ������������������������       �                      @                                   �?�����H�?             "@                                  �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?��
ц��?             :@                                 �?      �?             0@       ������������������������       �                     $@                                   �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@                                   �?z�G�z�?             9@                                   @K@      �?             0@        ������������������������       �                      @        ������������������������       �                     ,@                                   @J@�q�q�?             "@        ������������������������       �                     @                                  �U@      �?             @        ������������������������       �                     @        ������������������������       �                     @                +                    �?�z�G��?�             t@        !       (                   �r@��Q��?             D@       "       '                    �?     ��?             @@        #       &       
             �?�<ݚ�?             "@        $       %                     J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ,       O                   �b@�mTM�?�            �q@       -       D                    �?���[s�?�            �o@       .       3                   �c@���{h�?�            `l@       /       0                    `P@�6H�Z�?K            @]@       ������������������������       �        F             \@        1       2                    �P@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        4       ;                    �?�o�s(��?@            �[@        5       8                    �?�ݜ�?            �C@       6       7                 833@�g�y��?             ?@       ������������������������       �                     >@        ������������������������       �                     �?        9       :                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        <       =                    �?�J�T�?(            �Q@        ������������������������       �                     4@        >       C                    �?`'�J�?            �I@       ?       @       
             �?@9G��?            �H@        ������������������������       �                     6@        A       B                   �s@�>����?             ;@       ������������������������       �                     9@        ������������������������       �                      @        ������������������������       �                      @        E       F                    �?������?             ;@        ������������������������       �                     ,@        G       H                    �?��
ц��?
             *@        ������������������������       �                      @        I       L                    �?���|���?	             &@       J       K                 ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        M       N                     M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        P       S                   Po@�	j*D�?             :@        Q       R                   �e@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        T       W                     L@��S���?	             .@       U       V                   pg@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Y       �                    �?N����?�            �u@        Z       w                    �?X�Cc�?M             \@       [       b                    �?�d�����?6             S@        \       a                    �?j���� �?             1@       ]       `                   �a@�C��2(�?	             &@        ^       _                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        c       v                    �?�:�B��?+            �M@       d       s                   @e@"pc�
�?'            �K@       e       f                 ����?H%u��?%             I@        ������������������������       �                     2@        g       r                   s@     ��?             @@       h       m                   �b@�r����?             >@       i       j                   b@�nkK�?             7@       ������������������������       �                     1@        k       l                     M@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        n       o                    N@և���X�?             @        ������������������������       �                      @        p       q                   �n@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        t       u                   @`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        x       �                    �?X�<ݚ�?             B@       y       z                   �g@���@M^�?             ?@        ������������������������       �                     @        {       |                    @L@l��
I��?             ;@        ������������������������       �                     *@        }       �                   �?և���X�?	             ,@        ~                           �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@����X�?             @        �       �                   m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�K1T:�?�            @m@       �       �                    �?h�|׽?p             f@       �       �                   `[@4Jı@�?S            �_@        ������������������������       �                     >@        �       �                    �?��l��?C            @X@        �       �                 833�?��H�}�?             9@        ������������������������       �                     @        �       �                    �?�\��N��?             3@       �       �                 ����?���Q��?
             .@       �       �                   �`@      �?             (@        �       �                   �`@r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �a@r�q��?             @        ������������������������       �                     @        �       �                   0a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   m@������?4             R@       �       �                    �? >�֕�?            �A@        �       �                    b@�����H�?	             "@       ������������������������       �                     @        �       �                   `g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �? ��WV�?             :@        �       �                   �h@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                    �B@        ������������������������       �                     I@        �       �                    �?Ԫ2��?$            �L@       �       �                    `@r֛w���?             ?@       �       �                   @_@�q�q�?             8@       �       �                    �?z�G�z�?             4@        �       �                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �L@�t����?             1@        �       �                   �r@      �?              @       �       �                   �Y@      �?             @        ������������������������       �                     �?        �       �                    b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B�  ��1W-��?�<gTi��?���:*�??��W�?�������?�������?S֔5eM�?֔5eMY�?UUUUUU�?UUUUUU�?      �?                      �?�g�`�|�?L�Ϻ��?F]t�E�?]t�E�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?�؉�؉�?�;�;�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?������?�������?ffffff�?�������?      �?      �?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?              �?      �?        �_�_�?uPuP�?���p8�?����x<�?�9�K��?��gG�?�������?���?      �?        �������?�������?              �?      �?        �k߰��?J��yJ�?\��[���?�i�i�?��{���?�B!��?      �?                      �?      �?      �?      �?                      �?(�K=�?��V؜?      �?        �������?�?������?9/���?      �?        �Kh/��?h/�����?      �?                      �?      �?        B{	�%��?{	�%���?      �?        �؉�؉�?�;�;�?      �?        F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?                      �?vb'vb'�?;�;��?]t�E�?F]t�E�?      �?                      �?�?�������?�q�q�?�q�q�?      �?                      �?              �?DZ/`���?o)�'��?�m۶m��?%I�$I��?y�5���?Cy�5��?�������?ZZZZZZ�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?�pR���?�c+����?F]t�E�?/�袋.�?���Q��?)\���(�?              �?      �?      �?�?�������?d!Y�B�?�Mozӛ�?              �?UUUUUU�?�������?              �?      �?        ۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?      �?        �������?�������?              �?      �?                      �?r�q��?�q�q�?�s�9��?�c�1��?              �?Lh/����?h/�����?      �?        ۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?      �?                      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?�LɔLɴ?m�fm�f�?Cr��ѯ?�����?��b�X,�?O���t:�?              �?����?\���_�?
ףp=
�?{�G�z�?              �?�5��P�?y�5���?333333�?�������?      �?      �?�������?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�q�q�?�q�q�?�A�A�?��+��+�?�q�q�?�q�q�?              �?      �?      �?              �?      �?        ;�;��?O��N���?      �?      �?              �?      �?                      �?              �?              �?p�}��?$���>��?�B!��?���{��?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?�?<<<<<<�?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJA��2hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�6         b                 ����?�!���?�           ��@               C                    �?p���?�            Pw@                                  I@l-MIڼ�?�            0q@               	                    _@�����?             3@                                    I@ףp=
�?             $@                     
             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        
                            P@X�<ݚ�?             "@                                 @U@����X�?             @        ������������������������       �                     �?                                hff�?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               <                   �b@     G�?�             p@              7                   �t@@4և���?�            �m@              2                     P@�&xw���?�            @l@              %                    @L@��SПW�?�            �j@                                  �A@`���i��?j             f@                                   �?      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?                                  0n@Уp=
ע?_             d@       ������������������������       �        ;             Z@               $                   0d@�h����?$             L@              #       	             �?ܷ��?��?             =@                                 @[@d}h���?             ,@        ������������������������       �                      @                                    �I@�8��8��?
             (@       ������������������������       �                      @        !       "                    @J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             .@        ������������������������       �                     ;@        &       '                   �a@��-�=��?            �C@       ������������������������       �                     9@        (       1                     O@����X�?	             ,@       )       ,                    �L@���Q��?             $@        *       +                   �b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        -       .                   �i@���Q��?             @        ������������������������       �                      @        /       0                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        3       6                   Pc@�eP*L��?             &@       4       5                    ]@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        8       9       
             �?�q�q�?             (@       ������������������������       �                     @        :       ;                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        =       B                   �c@�<ݚ�?             2@        >       A                    �?z�G�z�?             @       ?       @                   0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        D       I                   P`@���c�H�?C            �X@        E       F                    �?`Ql�R�?             �G@       ������������������������       �                     F@        G       H                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       a                   �q@j���� �?#            �I@       K       T                    �?�p ��?            �D@       L       S                    �?8����?             7@       M       N                 ����?     ��?             0@        ������������������������       �                      @        O       P                   @d@      �?              @       ������������������������       �                     @        Q       R                   `g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        U       \                   �b@�<ݚ�?             2@        V       Y                    �?      �?             @        W       X                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       [                 lffֿ      �?             @        ������������������������       �                      @        ������������������������       �                      @        ]       `                   �_@�8��8��?             (@        ^       _                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     $@        c       �                   �b@�4�V�
�?�            �v@       d       w                    �?\-��p�?�             r@        e       r                    �?     x�?+             P@       f       m                   0`@��
ц��?            �C@       g       h                    \@z�G�z�?             4@        ������������������������       �                     &@        i       j                    �?X�<ݚ�?             "@        ������������������������       �                     @        k       l                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        n       q                   0b@�KM�]�?             3@       o       p                 033@�X�<ݺ?
             2@       ������������������������       �        	             1@        ������������������������       �                     �?        ������������������������       �                     �?        s       v                   Hw@HP�s��?             9@       t       u                   �X@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     �?        x       �                    �Q@0�֋���?�            @l@       y       �                    �?,N�_� �?�            �k@       z       �       
             �?HQ˄�ľ?�            @k@       {       �                    �?��R�x��?x            `g@        |                           �?�r����?	             .@        }       ~                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ����?�8��8��?             (@        ������������������������       �                     @        �       �                   @a@�����H�?             "@        ������������������������       �                     @        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��+��<�?o            �e@       �       �                 ����?�U���?P            �_@        �       �                   �`@�˹�m��?             C@       �       �                   `b@      �?             8@       �       �                 `ff�?      �?             0@        ������������������������       �                     @        �       �                   �r@�8��8��?             (@       ������������������������       �                     "@        �       �                     J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `c@      �?              @       �       �                    �?����X�?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �        9            @V@        �       �                   �_@��S�ۿ?            �F@        �       �                   @[@�q�q�?             @        ������������������������       �                     @        �       �                     M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����? ���J��?            �C@        �       �                   �q@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     :@        �       �                   P`@�n`���?             ?@        �       �                 ����?և���X�?             @        ������������������������       �                     �?        �       �                   �m@�q�q�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?      �?             8@        �       �                   `^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@P���Q�?             4@       ������������������������       �                     (@        �       �                    T@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �I@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @"` Y��?.            �Q@       �       �                    �?�d�����?#            �L@       �       �                    �?�Ra����?             F@       �       �                 ����?�+$�jP�?             ;@        �       �                   Pm@և���X�?             @       �       �                    �E@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   pe@P���Q�?
             4@       ������������������������       �        	             3@        ������������������������       �                     �?        ������������������������       �                     1@        �       �                    �?�θ�?	             *@       �       �                    �?և���X�?             @        ������������������������       �                     @        �       �                 ����?      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �B@d}h���?             ,@        ������������������������       �                     �?        �       �                    �N@8�Z$���?
             *@       ������������������������       �                     "@        �       �                   �c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  v��W�?E�q���?>N�� ��?�c����?���+�?�j����?^Cy�5�?Q^Cy��?�������?�������?�������?�������?              �?      �?                      �?r�q��?�q�q�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?              �?     `�?      �?n۶m۶�?�$I�$I�?v��\�(�?�8�1�s�?���o.��?��0�?F]t�E�?F]t�E�?      �?      �?      �?                      �?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?��=���?a���{�?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        }˷|˷�?�A�A�?      �?        �m۶m��?�$I�$I�?333333�?�������?�������?�������?              �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        t�E]t�?]t�E�?۶m۶m�?�$I�$I�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?9��8���?�q�q�?�������?�������?      �?      �?              �?      �?                      �?      �?        /�����?4և����?W�+�ɕ?}g���Q�?              �?UUUUUU�?UUUUUU�?      �?                      �?ZZZZZZ�?�������?dp>�c�?8��18�?8��Moz�?d!Y�B�?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?              �?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?ٞ u#�?J�w�"w�?�{a���?a����?      �?     ��?�;�;�?�؉�؉�?�������?�������?              �?�q�q�?r�q��?      �?        UUUUUU�?�������?      �?                      �?�k(���?(�����?��8��8�?�q�q�?      �?                      �?              �?{�G�z�?q=
ףp�?UUUUUU�?�������?      �?                      �?      �?        04��A�?�|٠ɗ�?���L�?h�`�|��?��p�?߅����?�и[�?��rD���?�?�������?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?w�qGܡ?�#�;��?��`0�?����|>�?^Cy�5�?��P^Cy�?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?              �?�?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?��-��-�?;�;��?�؉�؉�?              �?      �?                      �?�c�1��?�9�s��?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?      �?              �?      �?        �������?ffffff�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?              �?      �?              �?      �?        �V�H�?��RO�o�?Cy�5��?y�5���?]t�E]�?]t�E�?/�����?B{	�%��?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?        ffffff�?�������?      �?                      �?      �?        �؉�؉�?ى�؉��?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ojhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         �                    �?�#i����?�           ��@              -                    �?
j*D�?            z@               ,       	             �?L�];�?1            �Q@                                 �a@���e��?-            �P@                                   �?��
ц��?             :@              	                    i@
;&����?             7@                                  �R@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        
                          0r@����X�?             ,@                                  _@z�G�z�?	             $@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?              @                                  �?z�G�z�?             @        ������������������������       �                      @                                  @m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               !                    @G@��Q���?             D@                                  �b@      �?              @        ������������������������       �                     �?                                   �c@؇���X�?             @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        "       +                    �P@     ��?             @@       #       *                   @a@ 	��p�?             =@        $       )                   �`@"pc�
�?             &@       %       (                   �`@ףp=
�?             $@       &       '                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     @        ������������������������       �                     @        .       �                   hy@ )���?�            �u@       /       n       	             �?�����H�?�            `u@       0       1                 ����?�D?��7�?�            �s@        ������������������������       �        %            �P@        2       C                 ����? ��z)�?�            `o@        3       <                    �?b�2�tk�?             2@       4       ;                    �?      �?              @       5       :                    �?r�q��?             @       6       9                   p@      �?             @        7       8                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        =       B                   @d@z�G�z�?             $@       >       ?                 ����?�����H�?             "@        ������������������������       �                     @        @       A                   �\@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        D       ]       
             �?�ւ�?�?�             m@       E       \                    �R@�,���α?w            @h@       F       G                   h@��8����?v             h@        ������������������������       �        )             Q@        H       Q                    @G@`�c�г?M             _@        I       P                   @f@�r����?
             .@       J       K                    �?@4և���?	             ,@        ������������������������       �                     @        L       O                    �?      �?              @        M       N                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        R       Y                    c@бK/eh�?C            @[@       S       X                   @i@@䯦s#�?@            �Z@        T       U                    �?      �?             @        ������������������������       �                      @        V       W                   �h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        =            �Y@        Z       [                     O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ^       _                   pa@�(�Tw��?            �C@       ������������������������       �                     7@        `       m                    �?     ��?             0@       a       l                    �?X�Cc�?             ,@       b       k                    @�n_Y�K�?
             *@       c       d                   Pf@���!pc�?             &@        ������������������������       �                      @        e       j                    �?�����H�?             "@       f       g                 `ff�?      �?              @       ������������������������       �                     @        h       i                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        o       x                 833�?      �?             8@        p       q                    �?      �?              @        ������������������������       �                     �?        r       s                     C@����X�?             @        ������������������������       �                     �?        t       w                 ����?r�q��?             @       u       v                   `Y@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        y       �                    �?     ��?
             0@       z       �                   p`@z�G�z�?	             .@        {       �                    �?      �?             @       |                          d@���Q��?             @       }       ~                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                 033�D�E�?�            �s@        ������������������������       �                     @        �       �       	             �?���A�?�            �s@       �       �                 ���@Z,`��,�?�            �h@       �       �                    @O@�q���?�             h@       �       �                    �?����?q             d@       �       �                   �Q@$V�Ap�?c            �a@        ������������������������       �                      @        �       �                    �?��l��?b            �a@       �       �                   �b@T(y2��?U            �]@       �       �                    �? '��h�?P            @[@       �       �       
             �? �.�?Ƞ?.             N@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   pg@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        )             K@        �       �                    �?Hm_!'1�?"            �H@       �       �                    @K@�7��?            �C@       ������������������������       �                     ;@        �       �                 @33�?r�q��?	             (@       �       �                   pc@�����H�?             "@       ������������������������       �                     @        �       �                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?	             $@        ������������������������       �                     @        �       �                    @F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @k@�z�G��?             $@        ������������������������       �                     @        �       �                   Hq@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?���!pc�?             6@        ������������������������       �                     "@        �       �                 ����?��
ц��?	             *@       �       �                    �?�z�G��?             $@        �       �                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             2@        ������������������������       �                     @        �       �                   �l@      �?	             (@       ������������������������       �                     "@        ������������������������       �                     @        �       �                 833�?���@M^�?             ?@        �       �                    d@���Q��?             $@       �       �                    @P@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@����X�?             5@        �       �                    �?      �?             (@       �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �J@P����?O            �]@       ������������������������       �        2             S@        �       �                   pg@���N8�?             E@       �       �                   �?��Y��]�?            �D@       ������������������������       �                     >@        �       �                    @L@�C��2(�?             &@       ������������������������       �                     @        �       �                    �M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  �5�;���?%e��?��؉���?�؉�؉�?Zas �
�?SO�o�z�?>���>�?�>���?�;�;�?�؉�؉�?�Mozӛ�?Y�B��?9��8���?�q�q�?              �?      �?        �$I�$I�?�m۶m��?�������?�������?      �?      �?      �?                      �?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?      �?        �������?333333�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�{a���?������?F]t�E�?/�袋.�?�������?�������?UUUUUU�?�������?              �?      �?                      �?      �?                      �?      �?              �?        ��JVl�?á�=u2�?�q�q�?�q�q�?�1��X�?�J��?              �?G6q㓽?7>ّ�M�?�8��8��?9��8���?      �?      �?UUUUUU�?�������?      �?      �?      �?      �?      �?                      �?              �?              �?      �?        �������?�������?�q�q�?�q�q�?      �?        �������?UUUUUU�?              �?      �?                      �?�6���Ƴ?"9�A$��?���fy�?o�'�i��?�������?�����*�?              �?��RJ)��?��Zk���?�?�������?�$I�$I�?n۶m۶�?              �?      �?      �?      �?      �?              �?      �?                      �?      �?        ��A��.�?��]8��?�x+�R�?R����?      �?      �?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        � � �?�o��o��?              �?      �?      �?%I�$I��?�m۶m��?;�;��?ى�؉��?F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?              �?      �?      �?      �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?�������?�������?      �?      �?333333�?�������?      �?      �?      �?                      �?      �?                      �?              �?              �?      �?        q��;E�?=����?              �?gue*��?e*�kV��?T�r
^N�?�>4և��?UUUUU��?�������?���G��?���2��?�#T�ik�?��^���?              �?��O$���?f��k�?�F��F��?�5�5�?���]8��?�w� z|�?wwwwww�?�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        Y�Cc�?9/���?��[��[�?�A�A�?      �?        �������?UUUUUU�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ffffff�?333333�?      �?        �������?333333�?              �?      �?        F]t�E�?t�E]t�?      �?        �;�;�?�؉�؉�?ffffff�?333333�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        �s�9��?�c�1��?�������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?                      �?�V'u�?'u_[�?      �?        ��y��y�?�a�a�?8��18�?������?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��jhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKͅ�h��B@3         �       	             �?.��X~��?�           ��@              �       
             �?��%=�R�?j           X�@              D                    �?�7�%	�?           �z@               '                 ����?@g\:�?b            `d@               
                   @E@�99lMt�?.            �S@               	                    �J@r�q��?             (@                                  `_@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                  pc@���!pc�?(            �P@                                  �?@4և���?             E@                                  �?�?�|�?            �B@       ������������������������       �                     ?@                                   �?r�q��?             @                                  �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                ����?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                    @F@      �?             8@                                   �?      �?             (@        ������������������������       �                     �?                                   �?"pc�
�?             &@        ������������������������       �                     @                                   @C@�q�q�?             @        ������������������������       �                     �?                                   �D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        !       $                    �?      �?             (@        "       #                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        %       &                   f@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        (       C                    @�~6�]�?4            @U@       )       .                    �?����X�?)            �O@        *       -                    �?���Q��?             $@       +       ,                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        /       B                   �u@�T`�[k�?$            �J@       0       A                 033�?��x_F-�?"            �I@       1       4                    �?8��8���?              H@        2       3                     L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        5       >                   0e@�C��2(�?             F@       6       =                    �?@-�_ .�?            �B@       7       <                    �?HP�s��?             9@        8       ;                    c@"pc�
�?	             &@       9       :                    @O@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     (@        ?       @                    b@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        E       t                   0c@X�g�Y��?�            pp@       F       m                    �?���^���?�            �l@       G       l                    �?�g+��@�?�            �k@       H       S                    �?���Lͩ�?d            �b@        I       R                   b@�d�����?             3@       J       Q                   �`@     ��?             0@       K       P                   P`@      �?              @        L       M                    �?      �?             @        ������������������������       �                      @        N       O                    @H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        T       [                   �k@�	a�$a�?W            ``@        U       Z                    �? ������?+            �O@        V       Y                    �?P���Q�?             4@       W       X                    b@�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �E@        \       e                    \@�t����?,             Q@        ]       d                   �p@�n`���?             ?@        ^       _                    `@���Q��?             .@        ������������������������       �                     @        `       c                   �a@ףp=
�?             $@        a       b                   pm@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             0@        f       g                    �?@-�_ .�?            �B@       ������������������������       �                     ?@        h       k                   �`@�q�q�?             @        i       j                   p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        )             R@        n       o                   �Z@      �?              @        ������������������������       �                     �?        p       q                   `Z@؇���X�?             @       ������������������������       �                     @        r       s                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       ~                    d@:ɨ��?            �@@        v       }                 `ff@�q�q�?             (@       w       |                    �?z�G�z�?             $@       x       {                    �?�����H�?             "@        y       z                 033�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               �                    �?�����?             5@       �       �                   �r@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        �       �                   c@&� �N�?d             d@       �       �                   �`@4*T���?\            �b@        �       �                    �?8����?             G@       �       �                   @^@�IєX�?             A@        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     9@        ������������������������       �                     (@        �       �                   u@tt���A�?C            �Y@       �       �                 033�?z�G�z�?@            �W@       �       �                    �?,���i�?6            �T@        �       �                    �M@D�n�3�?             3@       �       �                 ����?և���X�?             ,@        ������������������������       �                     @        �       �                   �\@�q�q�?             "@        ������������������������       �                     @        �       �                    l@      �?             @        ������������������������       �                      @        �       �                   �_@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   Pt@�i�y�?(            �O@       �       �                   @[@0�z��?�?'             O@        �       �                    c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        $             M@        ������������������������       �                     �?        �       �                    �?�	j*D�?
             *@        ������������������������       �                     �?        �       �                    �?      �?	             (@       �       �                    �?�q�q�?             "@        �       �                    `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �s@r�q��?             (@       �       �                    �?�C��2(�?             &@       �       �                    �M@r�q��?             @        ������������������������       �                     @        �       �                    @P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   p@��<D�m�?a            `b@       �       �                     R@@�E�x�??            �X@       �       �                   �\@�a�O�?>            @X@        �       �                   �Z@      �?              @        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        7            @V@        ������������������������       �                     �?        �       �                 pff�?؇���X�?"            �H@       �       �                    �?�Ń��̧?             E@       ������������������������       �                     D@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                   Pb@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  ��� ���?���o���?O��v�&�?�0�ėl�?%�(f>�?��u&`��?K�m�
��?�ɀz��?5H�4H��?�o��o��?UUUUUU�?�������?�������?333333�?      �?                      �?              �?F]t�E�?t�E]t�?n۶m۶�?�$I�$I�?*�Y7�"�?к����?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        333333�?�������?      �?                      �?      �?      �?      �?      �?      �?        F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?r�q��?�q�q�?              �?      �?        �?999999�?�$I�$I�?�m۶m��?333333�?�������?�������?�������?      �?                      �?      �?        "5�x+��?���!5��?�?�������?�������?UUUUUU�?      �?      �?      �?                      �?F]t�E�?]t�E�?к����?S�n0E�?{�G�z�?q=
ףp�?F]t�E�?/�袋.�?�������?�������?              �?      �?              �?                      �?              �?�$I�$I�?�m۶m��?              �?      �?              �?              �?                      �?�x\�N�?�p�$��?���ϱ?ܯK*��?Nq��$�?���+c��?�K~��?�6�i�?y�5���?Cy�5��?      �?      �?      �?      �?      �?      �?              �?      �?      �?              �?      �?              �?                      �?              �?`�	)y��?T���0��?AA�?��}��}�?�������?ffffff�?�q�q�?��8��8�?              �?      �?                      �?              �?�?<<<<<<�?�c�1��?�9�s��?�������?333333�?      �?        �������?�������?UUUUUU�?�������?      �?                      �?              �?              �?к����?S�n0E�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?e�M6�d�?N6�d�M�?UUUUUU�?UUUUUU�?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?              �?                      �?              �?�a�a�?=��<���?�?�������?              �?      �?                      �?���2��?�l<�?�?w[��?�IA���?8��Moz�?d!Y�B�?�?�?�q�q�?9��8���?              �?      �?                      �?      �?        ����?��O ���?�������?�������?�����?8��18�?l(�����?(������?۶m۶m�?�$I�$I�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?      �?      �?              �?      �?                      �?      �?        �������?AA�?|���{�?�B!��?      �?      �?              �?      �?              �?                      �?;�;��?vb'vb'�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?        UUUUUU�?�������?F]t�E�?]t�E�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��S�r
�?և���X�?և���X�?9/���? tT����?����?      �?      �?      �?        �������?�������?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?��<��<�?�a�a�?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ9hExhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK酔h��B@:         �                    �?z��K���?�           ��@              [                   �c@�
�G�?           �{@              :                    �?d��G,�?�            �q@               /                    �?� ��1�?M            �^@              (       	             �?�'�`d�?>            �X@                                  �?�
��P�?5            @T@                                   �?      �?             <@                                   �?      �?             (@       	       
                   �_@      �?              @        ������������������������       �                     @                                  �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  0p@      �?             0@       ������������������������       �                     *@                                    M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�NW���?#            �J@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  `\@��<D�m�?            �H@                                  �R@�<ݚ�?             "@        ������������������������       �                     @                                   `P@      �?             @       ������������������������       �                      @        ������������������������       �                      @               '                   0h@�(\����?             D@                                    �?�}�+r��?
             3@        ������������������������       �                     "@        !       "                    �K@ףp=
�?             $@       ������������������������       �                     @        #       &                    �?�q�q�?             @       $       %                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        )       .                   �a@X�<ݚ�?	             2@       *       -                   �l@���!pc�?             &@       +       ,                   @_@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        0       9                    �R@      �?             8@       1       8                    �?���}<S�?             7@       2       7                    Y@؇���X�?
             ,@       3       6       	             �?�<ݚ�?             "@       4       5                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ;       J                   �e@X�Բ���?d            `d@        <       I                   �a@���>4��?             <@       =       D                    �?      �?             4@       >       C                 hff�?      �?             0@       ?       B                   @\@��S�ۿ?
             .@        @       A                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        E       H       	             �?      �?             @       F       G                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        K       P                    \@���?R            �`@        L       O                   �b@��<b���?             7@       M       N                    �N@ףp=
�?
             4@       ������������������������       �        	             2@        ������������������������       �                      @        ������������������������       �                     @        Q       R                     L@������?E             \@       ������������������������       �        1            �R@        S       T                    �L@�L���?            �B@        ������������������������       �                     �?        U       Z                 ����?�X�<ݺ?             B@       V       Y                    �M@�����?
             5@        W       X                   `p@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �        	             .@        \       �                 `ff@��T��g�?^            @c@       ]       l                    ]@̫���/�?Y            �a@        ^       k                    �?�	j*D�?             :@       _       d                   �h@��<b���?             7@        `       a                    �?      �?             @        ������������������������       �                      @        b       c                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        e       j                    �?�t����?
             1@       f       g                   `\@      �?	             0@       ������������������������       �                     ,@        h       i                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        m       ~                   �b@io8�?K             ]@       n       o                    �?X'"7��?E             [@       ������������������������       �        6            �U@        p       q                   �U@���N8�?             5@        ������������������������       �                     �?        r       }                    �?z�G�z�?             4@       s       z                    b@�����H�?             2@       t       u                    �?��S�ۿ?
             .@        ������������������������       �                     @        v       w                   Pe@ףp=
�?             $@        ������������������������       �                     @        x       y                   p`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        {       |                    l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               �                    �E@      �?              @        ������������������������       �                     �?        �       �                   0d@؇���X�?             @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        �       �                   �b@r�q��?�            `r@       �       �                    �?Ȱi�o��?�            Pp@       �       �                    �?�ւ�?�?�             m@        �       �                    �?j�q����?              I@       �       �                   @e@�ݜ�?            �C@       �       �       	             �?�8��8��?             B@       �       �                    �?h�����?             <@       �       �                   �]@�X�<ݺ?             2@       ������������������������       �                     (@        �       �                   P`@r�q��?             @        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �K@      �?              @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �R@�.ߴ#�?y            �f@       �       �                   �V@�ȉo(��?x            �f@        ������������������������       �                     �?        �       �                    �?�~
	�?w            �f@       �       �                   �h@ �&�eZ�?e             c@        ������������������������       �                     D@        �       �                    �? (��?K            @\@        �       �                   j@`'�J�?"            �I@        �       �                   �Y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��<b�ƥ?             G@        �       �                   �`@ףp=
�?             $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     B@        �       �                    �O@6uH���?)             O@       �       �                   ``@�1�`jg�?%            �K@       �       �                   �\@�8��8��?             B@        �       �                    �K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `@      �?             @@       �       �                   `a@(;L]n�?             >@        ������������������������       �        	             ,@        �       �                    �?      �?             0@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        �       �                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   �Z@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     <@        ������������������������       �                     �?        �       �                    �?���>4��?             <@        ������������������������       �                      @        �       �                 ����?      �?             4@        �       �                    �?      �?             @       �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?
             0@        ������������������������       �                      @        �       �                   @`@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�eP*L��?            �@@        �       �                    �?      �?             0@       �       �                   �l@r�q��?             (@       ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?������?	             1@        �       �                    @K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             (@        �       �                   �e@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �t�b�`     h�h)h,K ��h.��R�(KK�KK��hi�B�  K�ۚ��?�)|�� �?t�E]t�?]t�E�?D�{̒�?x��g��?������?������?'�l��&�?6�d�M6�?��ӭ�a�?������?      �?      �?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�x+�R�?萚`���?      �?      �?      �?                      �?և���X�?��S�r
�?�q�q�?9��8���?              �?      �?      �?              �?      �?        �������?333333�?(�����?�5��P�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?r�q��?�q�q�?t�E]t�?F]t�E�?      �?      �?              �?      �?                      �?      �?              �?      �?d!Y�B�?ӛ���7�?�$I�$I�?۶m۶m�?�q�q�?9��8���?      �?      �?      �?                      �?      �?                      �?              �?      �?        ��Ŗ��?kq�}�?I�$I�$�?n۶m۶�?      �?      �?      �?      �?�������?�?      �?      �?      �?                      �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?              �?��oS��?t��:W�?��,d!�?��Moz��?�������?�������?      �?                      �?              �?I�$I�$�?۶m۶m�?      �?        }���g�?L�Ϻ��?              �?��8��8�?�q�q�?=��<���?�a�a�?9��8���?�q�q�?      �?                      �?      �?              �?        �8+?!��?�S{��?Փ�ۥ��?Zas �
�?vb'vb'�?;�;��?��,d!�?��Moz��?      �?      �?      �?              �?      �?      �?                      �?<<<<<<�?�?      �?      �?      �?              �?      �?              �?      �?                      �?              �?|a���?GX�i��?Lh/����?B{	�%��?      �?        �a�a�?��y��y�?              �?�������?�������?�q�q�?�q�q�?�������?�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        UUUUUU�?�������?              �?      �?        UUUUUU�?�������?��;'�g�?e�� 3�?�6���Ƴ?"9�A$��?
ףp=
�?=
ףp=�?�i�i�?\��[���?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?�q�q�?��8��8�?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E]�?      �?                      �?XG��).�?�K�`m�?h�h��?�~��?      �?        >)7ͣ?�o��.��?�l�l�?�3��3��?              �?x�!���?H���?�?�������?�������?�������?      �?                      �?d!Y�B�?��7��M�?�������?�������?      �?      �?      �?                      �?              �?              �?��RJ)��?k���Zk�?�־a�?A��)A�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?      �?�?�������?              �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?      �?                      �?              �?      �?        n۶m۶�?I�$I�$�?      �?              �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?      �?              �?      �?        t�E]t�?]t�E�?      �?      �?�������?UUUUUU�?      �?        333333�?�������?      �?                      �?      �?        �?xxxxxx�?�������?�������?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ#9�*hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         �                    �?��;/M�?�           ��@              ;                   pa@~=�r�?           z@                                  �?���g<�?�            �q@                                  0m@�q�q�?             8@                                  �?���Q��?             .@        ������������������������       �                     @                                   @L@�q�q�?             "@       ������������������������       �                     @        	       
                   �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                ����?�����H�?             "@                                   �M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               ,                    �?`��F:u�?�            Pp@              +       
             �?�:�h���?�            �k@                                   �O@ �%�}��?y            �g@                                   E@ E��ۛ?^             b@                                   �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                   �?�|�l�?W             a@                                  \@����X�?F             \@                                  `_@ףp=
�?             $@       ������������������������       �                     @                                  �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        ?            �Y@        ������������������������       �                     8@        !       "                   �k@Du9iH��?            �E@        ������������������������       �                     3@        #       $                   @l@      �?             8@        ������������������������       �                      @        %       *                    �?���7�?             6@       &       )                   �Z@��S�ۿ?	             .@        '       (                 433�?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                    �@@        -       :       	             �?z�G�z�?             D@       .       /                    S@������?            �B@        ������������������������       �                     �?        0       7                   �r@�8��8��?             B@       1       2                   �]@Pa�	�?            �@@        ������������������������       �                     .@        3       6                 ����?�X�<ݺ?             2@        4       5                   @^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        8       9                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        <       k                   �`@�q�q�?V            �`@       =       `       
             �?��%��?0            �R@       >       W                   �p@`�Q��?#             I@       ?       R       	             �?4���C�?            �@@       @       M                    �J@X�Cc�?             <@       A       B                 ����?��.k���?             1@        ������������������������       �                     @        C       L                    �?X�Cc�?             ,@       D       E                    �C@�eP*L��?             &@        ������������������������       �                      @        F       G                    �?�q�q�?             "@        ������������������������       �                      @        H       I                    �?և���X�?             @        ������������������������       �                      @        J       K                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        N       O                    �O@�C��2(�?	             &@       ������������������������       �                     @        P       Q                   b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        S       V                    �J@z�G�z�?             @       T       U                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        X       _                   �e@�t����?             1@       Y       ^                    �?      �?
             0@       Z       [                    @G@@4և���?             ,@        ������������������������       �                     $@        \       ]                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        a       b                    �?      �?             8@        ������������������������       �                     (@        c       h                 033@      �?
             (@       d       e                   �k@      �?              @        ������������������������       �                      @        f       g                    b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        i       j                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        l       �                    �?д>��C�?&             M@        m       �                    �?      �?             @@       n                           �P@�q�q�?             8@       o       |                    �N@�ՙ/�?             5@       p       q                    �J@      �?
             0@        ������������������������       �                      @        r       y                    �?����X�?	             ,@       s       t                   �b@�����H�?             "@        ������������������������       �                     @        u       x                    �?�q�q�?             @       v       w       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        z       {       
             �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        }       ~                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	             �?$�q-�?             :@       �       �                   q@`2U0*��?             9@       ������������������������       �                     5@        �       �                    c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z��,i#�?�            �s@       �       �                 033��?�<��?�            @p@        ������������������������       �                     @        �       �       	             �?     ��?�             p@       �       �                    �?D>�Q�?c            �c@       �       �                   @E@����y7�?R            @_@        �       �                    �?��S���?             .@       �       �                   �X@���!pc�?             &@        ������������������������       �                     �?        �       �                    �?z�G�z�?             $@       �       �                    �M@      �?             @        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �O@���7�?G            �[@       �       �                    �?�K}��?A            �Y@       ������������������������       �        '             N@        �       �                    �?�Ń��̧?             E@        ������������������������       �                     *@        �       �                 433�?XB���?             =@       ������������������������       �                     :@        �       �                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @n@      �?              @        ������������������������       �                      @        �       �                   q@�q�q�?             @        ������������������������       �                     @        �       �                    `@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   hq@�g�y��?             ?@       �       �                   0c@������?             1@        ������������������������       �                     "@        �       �                   0d@      �?              @        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?d}h���?             ,@       ������������������������       �                     &@        ������������������������       �                     @        �       �                   @g@ �ׁsF�?B             Y@       ������������������������       �        A            �X@        ������������������������       �                     �?        �       �                 ����?�\��N��?!            �L@        �       �                   @`@R���Q�?             4@        �       �                   �]@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        �       �                 ����?����>�?            �B@       �       �                   �]@     ��?             @@        ������������������������       �                     $@        �       �                   �c@�eP*L��?             6@       �       �                   �X@      �?             0@        �       �                    �?�q�q�?             @       ������������������������       �                     @        �       �                   `b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 033�?z�G�z�?             $@       �       �                    �L@�����H�?             "@       ������������������������       �                     @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  �X�5��?�S�$e�?c�>ZMB�?gXp�l��?/<!W�³?z�����?�������?�������?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �q�q�?�q�q�?      �?      �?              �?      �?                      �?Ȥx�L��?�u�7[��?�*�*�?�F�F�?m�w6�;�?]AL� &�?����?�?�����?�q�q�?�q�q�?      �?                      �?~?�������?�$I�$I�?n۶m۶�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?w�qGܱ?qG�w��?              �?      �?      �?      �?        F]t�E�?�.�袋�?�?�������?UUUUUU�?�������?      �?                      �?              �?              �?              �?ffffff�?ffffff�?к����?��g�`��?      �?        UUUUUU�?UUUUUU�?|���?|���?              �?�q�q�?��8��8�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?}���g�?���L�?{�G�z�?��(\���?'�l��&�?m��&�l�?�m۶m��?%I�$I��?�������?�?              �?%I�$I��?�m۶m��?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?                      �?      �?        F]t�E�?]t�E�?              �?      �?      �?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?<<<<<<�?      �?      �?�$I�$I�?n۶m۶�?              �?      �?      �?      �?                      �?              �?      �?              �?      �?      �?              �?      �?      �?      �?              �?�������?UUUUUU�?              �?      �?              �?      �?              �?      �?        |a���?a���{�?      �?      �?UUUUUU�?UUUUUU�?�a�a�?�<��<��?      �?      �?              �?�$I�$I�?�m۶m��?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?333333�?�������?              �?      �?        �������?�������?      �?                      �?              �?              �?;�;��?�؉�؉�?{�G�z�?���Q��?              �?      �?      �?              �?      �?              �?        ��Sxǽ�?����?�����? �����?              �?     ��?      �?b'vb'v�?vb'vb'�?!�rh���?�~j�t��?�?�������?F]t�E�?t�E]t�?              �?�������?�������?      �?      �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?                      �?              �?�.�袋�?F]t�E�?�������?�?      �?        ��<��<�?�a�a�?      �?        GX�i���?�{a���?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�B!��?��{���?xxxxxx�?�?      �?              �?      �?              �?�������?�������?      �?                      �?۶m۶m�?I�$I�$�?              �?      �?        �G�z��?{�G�z�?      �?                      �?�5��P�?y�5���?333333�?333333�?�$I�$I�?۶m۶m�?      �?                      �?      �?        ���L�?�u�)�Y�?      �?      �?              �?]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�q�q�?�q�q�?      �?              �?      �?              �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJf/4'hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK煔h��B�9         z                    �?���-�g�?�           ��@                                  �?�u540��?�            0x@                                033�?D|U��@�?#            �P@               	                   �b@և���X�?             5@                                   �?"pc�
�?             &@        ������������������������       �                     �?                                  �l@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        
                           �?�z�G��?             $@                      	             �?���Q��?             @        ������������������������       �                      @                                  �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?��<b�ƥ?             G@                               ��� @�g�y��?             ?@                                   @K@�����H�?             "@                                  b@�q�q�?             @                                 `_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             6@        ������������������������       �                     .@               Y                 ����?���Q0�?�             t@              J                   �b@p��tKn�?�            �o@              -                    �?3e��?�            `m@              *                    �O@��AV���?d            �d@               '                   �?`#`��k�?^             c@       !       "       
             �?���=��?\            �b@       ������������������������       �        =             Z@        #       &                   c@��<b�ƥ?             G@        $       %                   �b@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     :@        (       )                   @a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        +       ,                   @t@����X�?             ,@       ������������������������       �                     $@        ������������������������       �                     @        .       C                    �?������?,             Q@       /       @                    �?�LQ�1	�?              G@       0       1                    �?$�q-�?            �C@        ������������������������       �                     ,@        2       5                   �^@H%u��?             9@        3       4                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        6       7                    _@�C��2(�?             6@        ������������������������       �                     @        8       9                    �I@�r����?             .@       ������������������������       �                     "@        :       ;                    `@�q�q�?             @        ������������������������       �                     �?        <       ?                   pf@z�G�z�?             @        =       >                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        A       B                   `\@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        D       E                     G@�eP*L��?             6@        ������������������������       �                     @        F       I                   �_@�t����?	             1@       G       H                     K@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        K       X                 @33�?�\��N��?             3@       L       U       	             �?��.k���?             1@       M       R                    �?�q�q�?             (@       N       O                    �?      �?              @        ������������������������       �                     @        P       Q                   Hq@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       T                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        V       W                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        Z       c                    �?�eP*L��?+            �P@        [       \                    �E@�t����?             1@        ������������������������       �                     �?        ]       ^                    �?      �?             0@       ������������������������       �                     (@        _       `                 ����?      �?             @        ������������������������       �                      @        a       b                   `T@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        d       m                    @K@~���L0�?            �H@        e       h                    �?r�q��?             8@       f       g                    @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        i       j                   �]@r�q��?             (@       ������������������������       �                      @        k       l                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        n       y                    �N@HP�s��?             9@       o       v                    c@�t����?             1@       p       q                    �M@@4և���?	             ,@       ������������������������       �                     @        r       s                   �]@؇���X�?             @        ������������������������       �                     @        t       u                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        w       x                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        {       �       	             �?h����?�            �u@       |       �                    �?�9����?�            �t@        }       �                   �`@N{�T6�?&            �K@        ~       �       
             �?��H�}�?             9@              �                   �b@      �?             2@       �       �                    �?�	j*D�?             *@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?r�q��?             >@       �       �                 ����?�����H�?             ;@       �       �                    @H@�S����?             3@        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �c@      �?             0@       ������������������������       �        	             ,@        �       �                   ps@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    `P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?��ś��?�            @q@       �       �                   Pb@      �?�             l@       �       �                    �?`�5���?            �g@        �       �                   �\@h�����?8             U@        �       �                   a@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                     Q@��pBI�?2            @R@       �       �                    �L@ ����?-            @P@        �       �                 ����?h�����?             <@        �       �                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                    �B@        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pl@�r�MȢ?G            �Z@       ������������������������       �        '             L@        �       �                   �[@`'�J�?             �I@        �       �                    �J@      �?             0@        ������������������������       �                     @        �       �                    Y@z�G�z�?             $@       ������������������������       �                     @        �       �                   �Z@�q�q�?             @       �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �A@        �       �                    �?���!pc�?            �@@       �       �                   �Z@�	j*D�?             :@        ������������������������       �                      @        �       �                    �?      �?             8@       �       �                 ����?d}h���?             ,@        ������������������������       �                     @        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                     M@�z�G��?             $@       ������������������������       �                     @        �       �                     P@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �I@؇���X�?             @       ������������������������       �                     @        �       �                    e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   p`@ s�n_Y�?             J@        �       �                   �b@և���X�?             5@       �       �                    `@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �l@z�G�z�?             $@        ������������������������       �                     @        �       �                   `m@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@`Jj��?             ?@       ������������������������       �                     9@        �       �                   @\@�q�q�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �^@      �?             0@        ������������������������       �                     @        �       �                 ����?�q�q�?             (@       ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                   d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  lk�w��?J��	.�?p�R,��? ��[���?�rv��?Xc"=P9�?۶m۶m�?�$I�$I�?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?        ffffff�?333333�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        d!Y�B�?��7��M�?�B!��?��{���?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?              �?              �?�����L�?�������?��`0�?����|>�?'�h��?�^��H��?��8���?7Āt,e�?@�?��?p�pŊ?�/��b��?O贁N{?      �?        ��7��M�?d!Y�B�?ffffff�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?xxxxxx�?�?��Moz��?Y�B��?�؉�؉�?;�;��?      �?        )\���(�?���Q��?UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        t�E]t�?]t�E�?              �?�������?�������?      �?      �?      �?                      �?      �?        y�5���?�5��P�?�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?              �?      �?              �?      �?      �?                      �?�������?�������?      �?                      �?      �?        ]t�E�?t�E]t�?<<<<<<�?�?              �?      �?      �?      �?              �?      �?      �?              �?      �?              �?      �?        ������?����>4�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?{�G�z�?q=
ףp�?�?<<<<<<�?�$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?����W��?ݏG*�?r'Gl���?$6�䈍�?pX���o�?�S�<%��?{�G�z�?
ףp=
�?      �?      �?vb'vb'�?;�;��?�������?333333�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?              �?      �?        UUUUUU�?�������?�q�q�?�q�q�?^Cy�5�?(������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        s��\;0�?R�g���?      �?      �?�d�hΚ?�ۤ��)�?�$I�$I�?�m۶m��?F]t�E�?]t�E�?              �?      �?        ����?���Ǐ�? �����? �����?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?              �?      �?      �?      �?                      �?�+J�#�?z����f�?              �?�?�������?      �?      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?t�E]t�?F]t�E�?;�;��?vb'vb'�?      �?              �?      �?۶m۶m�?I�$I�$�?              �?۶m۶m�?�$I�$I�?      �?                      �?333333�?ffffff�?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?�;�;�?۶m۶m�?�$I�$I�?F]t�E�?]t�E�?              �?      �?        �������?�������?      �?        333333�?�������?              �?      �?        �B!��?���{��?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJw�+hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         x                    �?�Fg�=��?�           ��@              i                    �?���!��?            {@              >                    �?�+$�jP�?�            �u@              	                    �?��ϻ�r�?�            `p@                                   �?��K2��?8            �W@                                   c@�g�y��?             ?@       ������������������������       �                     >@        ������������������������       �                     �?        ������������������������       �        )            �O@        
       7                    �?P����B�?u             e@                                 @[@z�G�z�?p             d@                                  �S@z�G�z�?             @        ������������������������       �                      @                                  �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               .                    �?�s�$$��?l            `c@                     	             �?ףp=
�?a            �a@                                   �?�����?,            �O@                                 �c@�O4R���?%            �J@                                 �c@`2U0*��?             9@       ������������������������       �                     8@        ������������������������       �                     �?        ������������������������       �                     <@                                  �l@      �?             $@        ������������������������       �                     @                                  �`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?               +                 033�?�s�c���?5            @S@                                  `X@�X�<ݺ?1             R@        ������������������������       �                     �?        !       *                    �?0z�(>��?0            �Q@       "       %                    �?���N8�?+            �O@        #       $                    �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        &       '                    @L@0�)AU��?'            �L@       ������������������������       �        !            �H@        (       )                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ,       -                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        /       0                 ����?�q�q�?             .@        ������������������������       �                     @        1       2                   �_@X�<ݚ�?             "@        ������������������������       �                      @        3       6                   �c@և���X�?             @       4       5                    �N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        8       9       	             �?      �?              @        ������������������������       �                     @        :       =                    �?���Q��?             @       ;       <                   e@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ?       P                   �`@4�<����?<            @V@        @       K                    �?�eP*L��?            �@@       A       F                   �h@      �?             4@        B       C                   �]@և���X�?             @        ������������������������       �                      @        D       E                   `_@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        G       J                    �?$�q-�?             *@        H       I                    Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        L       M                    `@�θ�?             *@       ������������������������       �                      @        N       O                    @E@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        Q       h                    �?���X�?%             L@       R       g                 ���@~���L0�?             �H@       S       \                    �?RB)��.�?            �E@       T       Y                    �?ܷ��?��?             =@        U       X                   pf@����X�?             @       V       W                    �G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        Z       [                   �b@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ]       ^                    @D@և���X�?             ,@        ������������������������       �                     @        _       f                   �r@���!pc�?             &@       `       a                 ����?      �?             @        ������������������������       �                      @        b       c                    �J@      �?             @        ������������������������       �                      @        d       e                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        j       k                   �O@j����?4            �T@        ������������������������       �                     <@        l       o                    �?D7�J��?            �K@       m       n                     N@$�q-�?             :@       ������������������������       �                     8@        ������������������������       �                      @        p       u       	             �?\-��p�?             =@       q       r                   �l@���}<S�?             7@       ������������������������       �                     (@        s       t                   �b@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        v       w                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        y       �                 hff�?,��4�?�            �r@        z       �                   �_@���|���?!            �K@        {       |                    �?�J�4�?             9@        ������������������������       �                     �?        }       ~       
             �?      �?             8@       ������������������������       �        	             0@               �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@��S���?             >@       �       �       
             �?�r����?
             .@       �       �                    �?@4և���?	             ,@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?z�G�z�?	             .@       �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�#-���?�            �n@       �       �                    �?@�qmNh�?s            `f@       �       �                    �?�̨�`<�?m            @e@       �       �                   �U@0��:�*�?[            �a@        ������������������������       �                      @        �       �                   p@Tri����?Z            �a@       �       �                   �e@�8��8��?>             X@       �       �                    �?���.�6�?;             W@        ������������������������       �                     &@        �       �                    �L@�>����?3            @T@       �       �                   P`@ �Cc}�?"             L@       �       �       
             �?     ��?             @@       �       �                    `@؇���X�?             <@       �       �                    @L@�C��2(�?             6@       �       �                    �?���N8�?             5@       �       �                    �?�}�+r��?             3@        �       �                   @Z@      �?              @        ������������������������       �                     @        �       �                    \@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   m@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     8@        ������������������������       �                     9@        �       �       
             �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?:	��ʵ�?            �F@       �       �                    @M@HP�s��?             9@       ������������������������       �                     2@        �       �                    �M@����X�?             @        ������������������������       �                     �?        �       �                   �`@r�q��?             @        �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �r@�z�G��?	             4@       �       �                   �p@�eP*L��?             &@       �       �       
             �?����X�?             @       �       �                    �K@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     ;@        �       �                   �t@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?����e��?,            �P@        �       �                    \@�nkK�?             7@        �       �                   @p@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                    �E@        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  �8�E$��?�c���?���M�&�?��Fd#��?/�����?B{	�%��?��6Ls�?qBJ�eD�?��Q�٨�?W�+�Ʌ?��{���?�B!��?      �?                      �?      �?        �a�a�?�y��y��?ffffff�?ffffff�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�����?�=���?�������?�������?=��<���?�a�a�?:�&oe�?�x+�R�?���Q��?{�G�z�?      �?                      �?      �?              �?      �?              �?�������?UUUUUU�?      �?                      �?�����?�cj`?��8��8�?�q�q�?              �?�ԓ�ۥ�?H���@��?��y��y�?�a�a�?UUUUUU�?UUUUUU�?              �?      �?        ��Gp�?p�}��?      �?              �?      �?              �?      �?              �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?      �?      �?      �?        �������?333333�?      �?      �?              �?      �?              �?        B�P�"�?|��^���?]t�E�?t�E]t�?      �?      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?              �?ى�؉��?�؉�؉�?      �?        �������?333333�?              �?      �?        ۶m۶m�?I�$I�$�?����>4�?������?S֔5eM�?���)k��?��=���?a���{�?�m۶m��?�$I�$I�?333333�?�������?              �?      �?              �?        �.�袋�?F]t�E�?      �?                      �?�$I�$I�?۶m۶m�?              �?F]t�E�?t�E]t�?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?        4u~�!��?f�@	o4�?              �?J��yJ�?k߰�k�?�؉�؉�?;�;��?      �?                      �?�{a���?a����?d!Y�B�?ӛ���7�?              �?F]t�E�?/�袋.�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ~��K~�?��:m��?F]t�E�?]t�E]�?{�G�z�?�z�G��?      �?              �?      �?              �?      �?      �?              �?      �?        �?�������?�������?�?n۶m۶�?�$I�$I�?�������?�������?              �?      �?              �?                      �?�������?�������?      �?      �?      �?                      �?              �?_�_�?�A�A�?�Fu��?I=W�l�?�?�������?�^���?H�>����?      �?        t�n���?�'Ni^�?UUUUUU�?UUUUUU�?Y�B��?���7���?              �?h/�����?�Kh/��?۶m۶m�?%I�$I��?      �?      �?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?�a�a�?��y��y�?(�����?�5��P�?      �?      �?              �?      �?      �?      �?      �?      �?                      �?              �?              �?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?        l�l��?��O��O�?{�G�z�?q=
ףp�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?333333�?ffffff�?t�E]t�?]t�E�?�$I�$I�?�m۶m��?�������?333333�?      �?                      �?              �?      �?                      �?              �?�q�q�?9��8���?              �?      �?        |���?�>����?d!Y�B�?�Mozӛ�?      �?      �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��+hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKӅ�h��B�4         \                 ����?�r,��?�           ��@              !                    �?�q�q�?�            pw@                                   �?r֛w���?J             _@                     	             �?�����	�?6            @U@                               833�?�˹�m��?0             S@       ������������������������       �        '            �O@                                   X@��
ц��?	             *@        ������������������������       �                     @        	       
                   �l@�q�q�?             "@       ������������������������       �                     @                                  0a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                  `n@�q�q�?             "@        ������������������������       �                     @                                  �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                ����?Hث3���?            �C@                                   �?      �?             (@        ������������������������       �                     @        ������������������������       �                     "@                                   `c@��}*_��?             ;@                                 �l@�eP*L��?
             6@        ������������������������       �                     @                                  �a@�q�q�?             2@        ������������������������       �                     @                                   �?؇���X�?             ,@       ������������������������       �                     "@                                  �p@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        "       Y                 ����?���w;�?�            `o@       #       4                   @E@dr����?�            �m@        $       3       	             �?X�<ݚ�?             2@       %       2                    `R@      �?             0@       &       1                    ^@�q�q�?             .@       '       (                    �J@�eP*L��?             &@        ������������������������       �                      @        )       0       
             �?�q�q�?             "@       *       /                    �?      �?              @       +       ,                     M@����X�?             @        ������������������������       �                     @        -       .                   �]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        5       H                    �?��`T.1�?�            �k@       6       E                   �f@@i�)ԙ�?y            �f@       7       @                   �? }�Я��?u            @f@       8       9                    �?�������?n            �d@       ������������������������       �        Z            �`@        :       ;                   �c@г�wY;�?             A@       ������������������������       �                     :@        <       =                   n@      �?              @        ������������������������       �                     @        >       ?                    @I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        A       D                    @M@�8��8��?             (@        B       C                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        F       G                   @b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        I       X       
             �?�q�q�?            �C@       J       S       	             �?|��?���?             ;@       K       R                   �b@     ��?             0@       L       Q                    �L@      �?	             $@       M       P                   �c@r�q��?             @        N       O                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        T       W                    @K@"pc�
�?             &@       U       V                   �g@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        Z       [                    �?�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        ]       �                    �?�?	���?�            pv@        ^                        033�?xk�2���?R            �_@       _       l                    �?�û��|�?+            @Q@        `       i       	             �?��a�n`�?             ?@       a       f                    �?H%u��?             9@       b       c                    @O@�}�+r��?
             3@       ������������������������       �                     (@        d       e                    @P@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        g       h                   �`@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        j       k                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        m       p                   �\@�\��N��?             C@        n       o                   �f@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        q       x                    �?�q�q�?             8@       r       s                    d@@4և���?             ,@       ������������������������       �                     "@        t       w                   �k@z�G�z�?             @        u       v                    e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        y       ~                    �?���Q��?             $@       z       }                 ����?X�<ݚ�?             "@       {       |                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �f@Riv����?'             M@       �       �                   pc@lGts��?&            �K@       �       �       	             �?���N8�?             E@       �       �                    @P@��Y��]�?            �D@       ������������������������       �                     B@        �       �       
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �c@�	j*D�?             *@        ������������������������       �                     �?        �       �                    @      �?
             (@        �       �                    o@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �R@�y��*�?�             m@       �       �                   �t@d����?�            �l@       �       �                    �?w��5o�?�            �j@        �       �                    �?      �?             @@       �       �                   @e@؇���X�?             <@       �       �                    �?�����H�?             ;@        ������������������������       �                     �?        �       �                 ����?$�q-�?             :@       �       �                    @F@8�Z$���?
             *@        ������������������������       �                      @        ������������������������       �        	             &@        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����@��?z            �f@       �       �                    �?*~k���?g            �b@       �       �                    �?r�q��?J             [@       �       �                   xt@��hJ,�?E            �Y@       �       �                   0c@�DÓ ��?D            @Y@       �       �                    �?�q��/��?B            �X@       �       �                   �U@����?-            @P@        ������������������������       �                     �?        �       �                    �L@     �?,             P@       �       �                   `_@@4և���?             E@       ������������������������       �                     6@        �       �                    �?R���Q�?             4@        ������������������������       �                      @        �       �                    �K@r�q��?             2@       �       �                   �a@�t����?             1@        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        �       �                    a@���Q��?             @       �       �                    l@      �?             @        ������������������������       �                      @        �       �                     I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                    �?r٣����?            �@@       �       �                 033�?�c�Α�?             =@        �       �                    @O@�eP*L��?             &@       �       �                    �F@����X�?             @        ������������������������       �                     �?        �       �                   �Y@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �J@r�q��?             2@        �       �                   �o@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                     @        �       �                   0p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    Z@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �E@        ������������������������       �                     >@        ������������������������       �                     1@        ������������������������       �                      @        �t�b�      h�h)h,K ��h.��R�(KK�KK��hi�B0  �292ȯ�?�f����?UUUUUU�?UUUUUU�?�B!��?���{��?�?{{{{{{�?^Cy�5�?��P^Cy�?              �?�؉�؉�?�;�;�?              �?UUUUUU�?UUUUUU�?      �?        �������?333333�?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �i�i�?��-��-�?      �?      �?      �?                      �?_B{	�%�?B{	�%��?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        333333�?�������?      �?                      �?      �?        ������?�핷$��?6�ф�?Tn�wpٻ?�q�q�?r�q��?      �?      �?UUUUUU�?UUUUUU�?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?      �?      �?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?      �?                      �?      �?              �?        �����?�����?��x��x�?��?�я~���?p�\��?(፦��?��k��x?      �?        �?�?      �?              �?      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?{	�%���?	�%����?      �?      �?      �?      �?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?/�袋.�?F]t�E�?333333�?�������?      �?                      �?      �?              �?        �������?�������?      �?                      �?X3��*�?*��M��?m6��f��?�d2�L&�?8��Moz�?��,d!�?�c�1��?�s�9��?)\���(�?���Q��?�5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�5��P�?y�5���?�$I�$I�?n۶m۶�?              �?      �?        �������?�������?n۶m۶�?�$I�$I�?      �?        �������?�������?      �?      �?              �?      �?              �?        �������?333333�?�q�q�?r�q��?UUUUUU�?�������?              �?      �?              �?                      �?	�=����?>�����?�־a�?�<%�S��?�a�a�?��y��y�?������?8��18�?              �?�������?�������?      �?                      �?      �?        ;�;��?vb'vb'�?      �?              �?      �?333333�?�������?      �?                      �?              �?      �?        GX�i��?�4�rO#�?�(�j�?�����a�?��n�?�?�-r�	�?      �?      �?�$I�$I�?۶m۶m�?�q�q�?�q�q�?      �?        ;�;��?�؉�؉�?;�;��?;�;��?      �?                      �?              �?      �?              �?        ��}kdu�?�C�rS��?�z=��?��^x/�?UUUUUU�?�������?�������?KKKKKK�?�~�X��?Q`ҩy��?և���X�?/����? �����?~�~��?      �?              �?     ��?�$I�$I�?n۶m۶�?              �?333333�?333333�?              �?UUUUUU�?�������?�?<<<<<<�?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?                      �?|���?>���>�?�{a���?5�rO#,�?]t�E�?t�E]t�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?                      �?UUUUUU�?�������?333333�?�������?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?              �?              �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���5hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B�5         �                    �?�Z���?�           ��@              q                    �?Ƞ����?n           �@              >                    �?�'�`d�?�            �r@               )                    �?      �?A             Z@              $                   �r@ގ�H��?.            �S@                                  �?���BK�?)            �Q@                     	             �?�99lMt�?            �C@              	                   pi@      �?             8@        ������������������������       �                     "@        
                          m@���Q��?             .@        ������������������������       �                     @                                   �?"pc�
�?             &@                                   o@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  Pm@��S���?             .@                                  �?�q�q�?             "@        ������������������������       �                     �?                                  �^@      �?              @        ������������������������       �                     @        ������������������������       �                      @                                   d@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �`@     ��?             @@       ������������������������       �                     5@                                  �a@�eP*L��?             &@                                  �o@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                !                   `c@r�q��?             @       ������������������������       �                     @        "       #                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        %       &                    �?      �?              @        ������������������������       �                     @        '       (                   xt@      �?             @        ������������������������       �                      @        ������������������������       �                      @        *       -                    b@� �	��?             9@        +       ,                   c@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        .       9                    `@�q�q�?             2@        /       6                    �?      �?              @       0       3       
             �?���Q��?             @        1       2       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       5                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       8                   �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        :       ;                   �c@z�G�z�?             $@       ������������������������       �                     @        <       =                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ?       T                    �?|�qh#��?~             h@        @       S                   �a@0B��D�?"            �M@       A       P                    �?�I� �?             G@       B       E                    �?���y4F�?             C@        C       D                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        F       G                    �?     ��?             @@        ������������������������       �                      @        H       K                    �E@      �?             8@        I       J                   �e@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        L       M                    @M@�IєX�?             1@       ������������������������       �                     *@        N       O                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        Q       R                     J@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        U       n                   �b@�iyw	
�?\            �`@       V       e                   @^@H*C�|F�?Y             `@        W       `                   �]@6uH���?)             O@       X       Y                    �? ��WV�?$             J@       ������������������������       �                     >@        Z       [                   �o@�C��2(�?             6@       ������������������������       �                     *@        \       ]                   �Y@�<ݚ�?             "@        ������������������������       �                     @        ^       _                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        a       b                    �?�z�G��?             $@       ������������������������       �                     @        c       d                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        f       m                    @J@0�,���?0            �P@        g       l                    �?�8��8��?             8@        h       i                    �H@�q�q�?             @        ������������������������       �                     �?        j       k                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                    �E@        o       p                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        r       �                   �?<��0�?�            @q@       s       �                   �b@88��M�?�            �j@       t       y                    �? �Jj�G�?G            �[@       u       x                    �?@�n���?B            �Y@        v       w                     Q@      �?             @@       ������������������������       �                     ?@        ������������������������       �                     �?        ������������������������       �        0            �Q@        z       {                   �c@؇���X�?             @        ������������������������       �                     @        |                           �?�q�q�?             @       }       ~                   n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @N@ȵHPS!�?C             Z@       �       �                    �?�$��y��?A            @X@       �       �       
             �?�(�Tw�?2            �S@       ������������������������       �                     �K@        �       �                    �?�nkK�?             7@        ������������������������       �                     @        �       �                   @[@�IєX�?             1@        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   �f@D�n�3�?             3@       �       �                   �c@և���X�?             ,@        ������������������������       �                     @        �       �                    �?�eP*L��?
             &@        ������������������������       �                     @        �       �                   n@      �?              @       �       �                   @i@      �?             @        ������������������������       �                     �?        �       �                   �j@���Q��?             @        ������������������������       �                     �?        �       �                   pf@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                     O@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @b@V{q֛w�?%             O@       �       �                    �?
;&����?             G@       �       �                   �U@ �o_��?             9@        ������������������������       �                     �?        �       �                   pa@      �?             8@        ������������������������       �                     &@        �       �                     K@��
ц��?             *@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��s����?             5@        ������������������������       �                      @        �       �                   0m@�KM�]�?
             3@       �       �                    �L@      �?             0@       ������������������������       �                     ,@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �\@     ��?
             0@        ������������������������       �                     @        ������������������������       �        	             *@        �       �                    �?���z��?j             d@       �       �                    �R@����W1�?M            @^@       �       �                   Pz@lZ�?��?L            @]@       �       �                   �c@ d�=��?J            @\@       �       �       
             �?`'�J�?C            �Y@       �       �                    �?p�C��?;            �V@       ������������������������       �        6            @T@        �       �                    �?z�G�z�?             $@       ������������������������       �                     @        �       �                 lffֿ�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@"pc�
�?             &@       ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   `d@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                   ``@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �U@��Q��?             D@        ������������������������       �        	             (@        �       �                     P@@4և���?             <@       �       �                    ]@ ��WV�?             :@        �       �                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�Bp  �H���x�?����C�?�#pi��??��-��?'�l��&�?6�d�M6�?      �?      �?��td�@�?���M���?$Zas �?��RO�o�?�o��o��?5H�4H��?      �?      �?              �?�������?333333�?      �?        F]t�E�?/�袋.�?      �?      �?      �?                      �?              �?�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?UUUUUU�?              �?      �?              �?      �?              �?]t�E�?t�E]t�?�������?�������?      �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?�Q����?)\���(�?�$I�$I�?�m۶m��?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?333333�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�n�տ?=RBN�?��}ylE�?�A�I��?Nozӛ��?Y�B���?(������?6��P^C�?�������?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?�$I�$I�?�m۶m��?              �?      �?        �?�?              �?      �?      �?              �?      �?              �?      �?              �?      �?                      �?*g��1�?����?�!oȫ?�7�yC�?��RJ)��?k���Zk�?;�;��?O��N���?              �?F]t�E�?]t�E�?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?ffffff�?              �?      �?      �?      �?                      �?g��1��?Ez�rv�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?              �?�������?333333�?              �?      �?        4J��?�?0�̵�?+J�#��?����f��?k߰�k�?��)A��?\mMw��?��,�?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ��N��N�?�؉�؉�?����?W?���?p��o���?�A�A�?      �?        �Mozӛ�?d!Y�B�?      �?        �?�?      �?      �?              �?      �?              �?        l(�����?(������?۶m۶m�?�$I�$I�?              �?t�E]t�?]t�E�?      �?              �?      �?      �?      �?              �?333333�?�������?      �?              �?      �?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?        B!��?�{����?�Mozӛ�?Y�B��?
ףp=
�?�Q����?              �?      �?      �?      �?        �;�;�?�؉�؉�?      �?                      �?�a�a�?z��y���?      �?        (�����?�k(���?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        ��6��?\|r��?���|���?��eP*L�?^�^�?=�C=�C�?x�!���?���	��?�?�������?h�h��?��K��K�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?        F]t�E�?]t�E]�?      �?                      �?      �?      �?              �?      �?              �?        �������?ffffff�?              �?n۶m۶�?�$I�$I�?O��N���?;�;��?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJRܯ[hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�6         �                    �?���:���?�           ��@              m                   �b@h����)�?           0y@                                 Pf@��̃Z�?�            u@                                  `f@ ���J��?E            @]@                                  �?�Ru߬Α?C            �\@                                   @K@Pa�	�?            �@@               
                    �?ףp=
�?             $@               	                    @J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �        0            @T@                                    O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               ,                    �?��#:���?�            �k@               #                   xp@�z�6�?.             O@                                  �?r�q��?$             H@                                   @N@      �?              @        ������������������������       �                      @                                   `P@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @                                  0`@ףp=
�?             D@       ������������������������       �                     6@                                  p`@�<ݚ�?             2@        ������������������������       �                     �?                                   `@@�0�!��?             1@        ������������������������       �                     @               "                   0a@�z�G��?             $@                !                   Pb@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        $       )                   Hq@X�Cc�?
             ,@        %       (       	             �?z�G�z�?             @       &       '                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        *       +                   �Y@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        -       F                    `@�v,D�?n            �c@        .       E                    �?�%^�?            �E@       /       D       
             �?��P���?            �D@       0       3                 ����?�I�w�"�?             C@        1       2                 ����?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        4       =                    �?"pc�
�?            �@@       5       6                    �?������?             1@        ������������������������       �                     @        7       <                    �J@����X�?
             ,@        8       ;                     @�q�q�?             @       9       :                    @G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        >       C                   P`@      �?             0@        ?       B                   `_@���Q��?             @       @       A                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        G       H                   �f@���}<S�?O            �\@        ������������������������       �                     �?        I       ^                   pn@�˹�m��?N            �\@        J       ]       	             �?r�q��?             E@       K       P                    �?�p ��?            �D@        L       M                    �?      �?              @       ������������������������       �                     @        N       O                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        Q       V                 `ff�?�C��2(�?            �@@        R       U                   `m@���Q��?             @       S       T                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        W       \                 ����?h�����?             <@        X       Y                    �?r�q��?             @        ������������������������       �                     @        Z       [                   @\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     �?        _       h                    �?������?0             R@       `       g                   ``@ ����?+            @P@        a       f                 ����?�C��2(�?             &@       b       e                    �?z�G�z�?             @       c       d                    �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        #             K@        i       l                   @^@؇���X�?             @       j       k                   �Z@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        n                           �?�'�=z��?,            �P@       o       x                   �n@\�Uo��?             C@       p       w       	             �?�+e�X�?             9@       q       r                   �Q@�z�G��?             4@        ������������������������       �                     @        s       t       
             �?@�0�!��?             1@        ������������������������       �                     �?        u       v                    @      �?             0@       ������������������������       �        
             ,@        ������������������������       �                      @        ������������������������       �                     @        y       z       
             �?�	j*D�?	             *@        ������������������������       �                     @        {       ~                   �p@�q�q�?             @       |       }                     E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   c@��X��?             <@        ������������������������       �                      @        �       �                    q@R�}e�.�?             :@       ������������������������       �        	             ,@        �       �                 @33�?�q�q�?             (@        ������������������������       �                     @        �       �                   y@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @E@��>K��?�            �t@        �       �                 hff�?      �?             B@       �       �                    �?j���� �?             1@       �       �                 ����?�<ݚ�?             "@       �       �                    �P@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�KM�]�?
             3@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        �       �                    �?΂.o�?�            pr@       �       �                   �?�p8[(��?�             n@       �       �                    @M@��e�_�?u            �g@       �       �       	             �?�C��2(�?j             f@       �       �                   0n@      �?7             X@       ������������������������       �        &             O@        �       �                 ����?l��\��?             A@       �       �                    �? �Cc}�?             <@       �       �                    o@$�q-�?             :@        ������������������������       �                      @        ������������������������       �                     8@        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        3             T@        �       �                    �?8�Z$���?             *@       ������������������������       �                     "@        �       �                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �^@ s�n_Y�?              J@        ������������������������       �                     @        �       �                    �?ZՏ�m|�?            �H@       �       �                    �?�����H�?             B@        ������������������������       �                     $@        �       �       	             �?8�Z$���?             :@       �       �                    �?$�q-�?	             *@       ������������������������       �                     $@        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     L@�θ�?             *@       ������������������������       �                      @        �       �                   p`@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�	j*D�?             *@       �       �                    @"pc�
�?             &@       �       �                   �^@ףp=
�?             $@        ������������������������       �                     @        �       �                   pi@      �?             @        ������������������������       �                      @        �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?J��D��?)             K@       �       �                    �? >�֕�?            �A@        ������������������������       �                     0@        �       �                   �c@�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @        �       �                    �?���y4F�?             3@        �       �                   �a@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    @K@�r����?             .@        �       �                    �?����X�?             @       �       �                    @F@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   `e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  !��Q��?p��1W-�?�f��?�<�Ef��?���X�?���|�?�A�A�?��-��-�?p�}��?���#��?|���?|���?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?�S�<%��?k߰��?�Zk����?J)��RJ�?UUUUUU�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?�q�q�?9��8���?      �?        �������?ZZZZZZ�?              �?333333�?ffffff�?333333�?�������?      �?                      �?              �?�m۶m��?%I�$I��?�������?�������?      �?      �?              �?      �?              �?        �q�q�?�q�q�?      �?                      �?�ґ=�?~W��0��?�}A_�?�}A_��?�����?������?�5��P�?����k�?333333�?�������?              �?      �?        F]t�E�?/�袋.�?�?xxxxxx�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?�������?333333�?      �?      �?      �?                      �?      �?                      �?              �?      �?        d!Y�B�?ӛ���7�?      �?        ^Cy�5�?��P^Cy�?UUUUUU�?�������?��+Q��?Q��+Q�?      �?      �?              �?      �?      �?      �?                      �?F]t�E�?]t�E�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �q�q�?�q�q�? �����? �����?F]t�E�?]t�E�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?|���?|��|�?�5��P^�?6��P^C�?R���Q�?���Q��?ffffff�?333333�?              �?ZZZZZZ�?�������?              �?      �?      �?      �?                      �?      �?        ;�;��?vb'vb'�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        %I�$I��?n۶m۶�?      �?        �;�;�?'vb'vb�?              �?�������?�������?              �?      �?      �?      �?                      �?.��3�?F�\��3�?      �?      �?ZZZZZZ�?�������?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?(�����?�k(���?UUUUUU�?UUUUUU�?              �?      �?                      �?�o�U�k�?o��P%��?�!��!��?�����?t���G'�?p����?t�E]t�?t�E]t�?      �?      �?      �?        ------�?�������?%I�$I��?۶m۶m�?�؉�؉�?;�;��?              �?      �?              �?      �?              �?      �?              �?              �?        ;�;��?;�;��?      �?              �?      �?      �?                      �?�;�;�?;�;��?              �?�>4և��?9/����?�q�q�?�q�q�?      �?        ;�;��?;�;��?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ى�؉��?�؉�؉�?      �?        �������?333333�?              �?      �?        vb'vb'�?;�;��?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?      �?              �?      �?              �?      �?                      �?              �?�^B{	��?_B{	�%�?��+��+�?�A�A�?      �?        �k(���?(�����?      �?                      �?(������?6��P^C�?      �?      �?      �?                      �?�?�������?�$I�$I�?�m۶m��?�������?�������?              �?      �?              �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ[P!hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK酔h��B@:         t                 ����?�$���?�           ��@              k                    �?���3�g�?�             w@              B                    @L@TI�M���?�            v@              ;                    �?      �?�             p@                                  �?��<b���?�            �l@                                  @G@�:�]��?b             c@        ������������������������       �        ,            �P@                                  @[@\-��p�?6            �U@        	                           i@r�q��?             @       
              	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   �? wVX(6�?3            @T@                               ����?`����֜?,            �Q@                                  �?��v$���?&            �N@       ������������������������       �        !             J@                                  `f@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@                                  @a@�eP*L��?             &@                               ����?����X�?             @                     	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               .                    �?�J���?/            @S@                                  �?�P�*�?"             O@        ������������������������       �                     4@                '                    �?؇���X�?             E@        !       "                   e@R���Q�?             4@       ������������������������       �                     &@        #       $                    �?�q�q�?             "@        ������������������������       �                      @        %       &                   0j@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        (       -                   @b@��2(&�?             6@       )       ,                    @F@�����?             5@        *       +                   �[@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     �?        /       8                    �?z�G�z�?             .@       0       1                   �`@r�q��?
             (@        ������������������������       �                     @        2       3                    �?�q�q�?             @        ������������������������       �                     �?        4       7                   �a@z�G�z�?             @        5       6                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        9       :                    @G@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        <       A                    �?��
ц��?             :@       =       >                    �z�G�z�?             .@        ������������������������       �                      @        ?       @                    @E@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     &@        C       T                    �?�U�!��?A            @X@        D       Q                    �?�������?             F@        E       P                   �b@�ՙ/�?             5@       F       G                    �?     ��?             0@        ������������������������       �                     �?        H       O       	             �?�r����?
             .@       I       J                   �a@@4և���?	             ,@       ������������������������       �                     $@        K       N                    �?      �?             @       L       M                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        R       S                   Pa@�nkK�?             7@       ������������������������       �                     6@        ������������������������       �                     �?        U       V                    �?�c�����?&            �J@       ������������������������       �                     ?@        W       j                    �P@8�A�0��?             6@       X       e                   �c@      �?             2@       Y       d                    �?z�G�z�?
             $@       Z       a                    �?����X�?             @       [       \                    �?z�G�z�?             @        ������������������������       �                      @        ]       ^                   �^@�q�q�?             @        ������������������������       �                     �?        _       `                   `X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        b       c                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        f       g                   �d@      �?              @       ������������������������       �                     @        h       i                   `@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        l       s                    �?ҳ�wY;�?	             1@       m       r                    �?���Q��?             .@       n       o                   `c@ףp=
�?             $@       ������������������������       �                      @        p       q                   p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        u       �                    �?d}h���?�            �v@        v       �                    �J@6C�z��?M            �\@        w       �                    b@�������?             A@       x       �                 ����?؇���X�?             <@       y       �                    �?����X�?             ,@       z                          �d@�θ�?             *@       {       |                 pff�?ףp=
�?	             $@       ������������������������       �                      @        }       ~                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `P@�z�Ga�?3             T@       �       �                    �?d,���O�?&            �I@       �       �                    �?R���Q�?             D@       �       �                    �?�#-���?            �A@       ������������������������       �                     8@        �       �                   Xr@���!pc�?	             &@       ������������������������       �                     @        �       �                    b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   0c@���Q��?             @       �       �                   �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �L@���|���?
             &@        ������������������������       �                     @        �       �                   �e@�q�q�?             @       �       �                   �b@      �?             @        ������������������������       �                     �?        �       �                    j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �R@����"�?             =@       �       �                    �?
j*D>�?             :@        ������������������������       �                     &@        �       �                   �b@������?             .@       �       �                    �?8�Z$���?             *@        �       �                   �n@����X�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �R@h�N?���?�            @o@       �       �                    �?�}#���?�             o@        �       �                   P`@���y4F�?             C@        �       �                   �\@      �?             $@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �`@ �Cc}�?             <@       ������������������������       �                     6@        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   @^@8�W���?�            `j@        �       �                   Hs@�:�B��?"            �M@       �       �                    �?؇���X�?              L@       �       �                   �U@ףp=
�?             I@        ������������������������       �                     �?        �       �                 033�?Hm_!'1�?            �H@        ������������������������       �        	             0@        �       �                    �?<���D�?            �@@       �       �                    @L@@4և���?             <@       ������������������������       �        
             2@        �       �                    �M@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @       �       �                   �n@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �i@pe�D�ϣ?a             c@        �       �                    �?`�q�0ܴ?            �G@       �       �                    �? �#�Ѵ�?            �E@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@��Y��]�?            �D@       �       �                    �?���7�?             6@       ������������������������       �        	             .@        �       �                   �Y@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             3@        ������������������������       �                     @        �       �                    @M@@��!�Q�?D            @Z@       ������������������������       �        (            @P@        �       �                    c@�(\����?             D@       ������������������������       �                     C@        �       �                   `o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B�  �E$�~V�?�����?�UҨ�\�?iT[��F�?� �����?����RN�?      �?      �?��,d!�?��Moz��?}}}}}}�?�?      �?        a����?�{a���?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?k~X�<�?�<ݚ�?�������?�A�A�?.�u�y�?;ڼOqɐ?      �?        �q�q�?�q�q�?      �?                      �?      �?        ]t�E�?t�E]t�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?����15�?qV~B���?�RJ)���?�Zk����?              �?۶m۶m�?�$I�$I�?333333�?333333�?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?        ��.���?t�E]t�?=��<���?�a�a�?333333�?�������?              �?      �?              �?                      �?�������?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?�;�;�?�������?�������?              �?�؉�؉�?;�;��?              �?      �?                      �?���:*�? tT����?/�袋.�?t�E]t�?�a�a�?�<��<��?      �?      �?      �?        �?�������?�$I�$I�?n۶m۶�?              �?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        d!Y�B�?�Mozӛ�?              �?      �?        �V�9�&�?:�&oe�?      �?        /�袋.�?颋.���?      �?      �?�������?�������?�m۶m��?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?�������?333333�?�������?�������?              �?      �?      �?      �?                      �?      �?                      �?۶m۶m�?I�$I�$�?��Gp�?~��G�?�������?�������?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?ى�؉��?�؉�؉�?�������?�������?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?�������?              �?      �?        �������?�������?PPPPPP�?�������?333333�?333333�?_�_�?�A�A�?              �?t�E]t�?F]t�E�?              �?333333�?�������?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?	�=����?�i��F�?b'vb'v�?;�;��?      �?        �?wwwwww�?;�;��?;�;��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?              �?        �I+��?�v��/�?4u~�!��?Y1P�M�?(������?6��P^C�?      �?      �?              �?�������?UUUUUU�?      �?                      �?۶m۶m�?%I�$I��?              �?      �?      �?      �?                      �?��H����?Cs;�G�?�pR���?�c+����?�$I�$I�?۶m۶m�?�������?�������?      �?        9/���?Y�Cc�?              �?|���?|���?�$I�$I�?n۶m۶�?              �?�������?�������?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?^Cy�5�?�5��P^�?W�+�ɥ?��F}g��?�}A_Ч?�/����?      �?      �?              �?      �?        ������?8��18�?F]t�E�?�.�袋�?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?8�8��? �����?              �?�������?333333�?              �?      �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��,@hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKÅ�h��B�0         l                    �?j8je3�?�           ��@              #                    �?B�a���?           py@               "       	             �?�������?'             N@                                  a@x�K��?!            �I@                                 �[@      �?             8@                                  �e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        	                           �?�d�����?             3@       
                          0n@z�G�z�?             .@        ������������������������       �                      @                                   �?և���X�?             @                                  @H@���Q��?             @        ������������������������       �                     �?                                   �?      �?             @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                    M@      �?             @        ������������������������       �                      @        ������������������������       �                      @               !                    �?�+$�jP�?             ;@                                   `P@X�Cc�?	             ,@                                 �x@"pc�
�?             &@       ������������������������       �                      @                                   @O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     "@        $       _                    �?������?�            �u@       %       @                    �?@��3�2�?�            �q@        &       -                    @F@8�Z$���?5            �S@        '       ,                    @X�<ݚ�?             "@       (       +                    �?և���X�?             @        )       *                     C@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        .       /                   `k@ ���g=�?-            @Q@        ������������������������       �                     ?@        0       ;       	             �?���y4F�?             C@       1       :                   �`@���}<S�?             7@        2       9                    �?�<ݚ�?             "@       3       4                    @L@����X�?             @        ������������������������       �                     @        5       6                     N@�q�q�?             @        ������������������������       �                     �?        7       8                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             ,@        <       ?                   `n@���Q��?             .@       =       >                     J@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        A       N                    �?����?�            @i@        B       G                    �?H%u��?             9@        C       D                    �?���Q��?             @        ������������������������       �                     �?        E       F                    �L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        H       M                   �U@P���Q�?             4@        I       L                    @K@      �?              @        J       K                    W@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        O       P                    @K@����7�?u             f@        ������������������������       �        7            @U@        Q       ^                   �a@��<b�ƥ?>             W@       R       ]                    �?�&=�w��?%            �J@       S       V                    �?@-�_ .�?            �B@        T       U                   a@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        W       \                   �[@�g�y��?             ?@        X       [                    �?r�q��?             @        Y       Z                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@        ������������������������       �                     0@        ������������������������       �                    �C@        `       i                   �b@h��Q(�?*            �P@       a       b                 ����?      �?             H@       ������������������������       �                     9@        c       h                    �?�LQ�1	�?             7@        d       g                    �?      �?             @       e       f                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             3@        j       k                   8p@D�n�3�?             3@       ������������������������       �                     &@        ������������������������       �                      @        m       �                    �? ��?�?�            pt@       n       �                    �?6&�����?�            Pp@       o       �                   h@$�q-�?y            �f@       p       �                 ���@�O2�J�?w             f@       q       �                   �a@��-��ĳ?v            �e@       r       {                   �a@PL��V�?b            �b@        s       t                    �?�nkK�?             G@        ������������������������       �                     5@        u       v                    @L@HP�s��?             9@       ������������������������       �                     2@        w       x                 @33�?����X�?             @        ������������������������       �                      @        y       z                   p`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        |       }                   �`@�K}��?C            �Y@       ������������������������       �        0             S@        ~       �                   �`@ ��WV�?             :@               �                 ����?�q�q�?             @        ������������������������       �                     �?        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?8�Z$���?             :@       �       �                   �_@�����?             5@        �       �                    ^@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        �       �                    �P@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?v�_���?1            �S@       �       �                    �?�θ�?(            @P@        �       �                    �M@d��0u��?             >@       �       �                   �_@�	j*D�?             :@       �       �                    @J@�n_Y�K�?
             *@       �       �                    �?      �?             $@       �       �                   0l@����X�?             @        ������������������������       �                     @        �       �                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        �       �                   �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `P@(N:!���?            �A@       �       �                   �_@      �?             @@        �       �                   �[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     <@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    `@؇���X�?	             ,@       ������������������������       �                     (@        ������������������������       �                      @        �       �                   Pd@�{r٣��?$            �P@       �       �                    c@`��}3��?            �J@       �       �       
             �?�*/�8V�?            �G@       �       �                    �N@��-�=��?            �C@       �       �                    �?PN��T'�?             ;@        ������������������������       �                      @        �       �                   �b@HP�s��?             9@       �       �                   �_@ �q�q�?             8@        �       �                   q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             2@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        �       �                    @M@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KK�KK��hi�B0  ���Y��?t�S��?�s�ө��?��UH�?�������?�������?�?ssssss�?      �?      �?�������?�������?              �?      �?        Cy�5��?y�5���?�������?�������?      �?        �$I�$I�?۶m۶m�?�������?333333�?              �?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?      �?              �?      �?              �?      �?        B{	�%��?/�����?�m۶m��?%I�$I��?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ��X�޶?��\&$�?_�_��?���?;�;��?;�;��?�q�q�?r�q��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?                      �?ہ�v`��?��(�3J�?              �?(������?6��P^C�?d!Y�B�?ӛ���7�?�q�q�?9��8���?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?�������?333333�?      �?      �?              �?      �?                      �?z��~�X�?|#
L:5�?���Q��?)\���(�?�������?333333�?      �?              �?      �?              �?      �?        �������?ffffff�?      �?      �?      �?      �?      �?                      �?              �?              �?��F($�?��^o��?              �?d!Y�B�?��7��M�?�x+�R�?tHM0���?к����?S�n0E�?UUUUUU�?�������?              �?      �?        �B!��?��{���?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?              �?              �?z�rv��?�Wc"=P�?      �?      �?              �?Y�B��?��Moz��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?l(�����?(������?      �?                      �?߅���]�?���]8��?�<ZT"��?���v�?�؉�؉�?;�;��?�v�,1�?k��2�?�f��o��?/�I���?�u�)�Y�?L�Ϻ��?�Mozӛ�?d!Y�B�?      �?        q=
ףp�?{�G�z�?      �?        �m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?        �������?�?      �?        O��N���?;�;��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        ;�;��?;�;��?=��<���?�a�a�?UUUUUU�?UUUUUU�?      �?                      �?      �?        333333�?�������?      �?                      �?              �?�������?�������?      �?                      �? *�3�?���M���?ى�؉��?�؉�؉�?DDDDDD�?wwwwww�?vb'vb'�?;�;��?ى�؉��?;�;��?      �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?      �?              �?      �?        |�W|�W�?�A�A�?      �?      �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        |���?��|��?M0��>��?�琚`��?AL� &W�?�٨�l��?�A�A�?}˷|˷�?h/�����?&���^B�?      �?        {�G�z�?q=
ףp�?UUUUUU�?�������?UUUUUU�?�������?              �?      �?                      �?      �?                      �?      �?        �������?UUUUUU�?              �?      �?        �؉�؉�?;�;��?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��PhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKх�h��B@4         H                   �`@����?�           ��@               5                    �?���N8�?�             u@                                  �?������?�            0p@                                   �?D�n�3�?             3@              
                    �H@     ��?             0@                                   �G@      �?             @        ������������������������       �                     �?               	                   �k@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �a@r�q��?             (@       ������������������������       �                     "@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               4                   �z@��*;�?�             n@              3                    �R@�����?�            �m@                                  @L@��Uu ְ?�            `m@        ������������������������       �        A             Z@               ,                    �?�-�[�?N            ``@              +                 ����?P���Q�?I             ^@              $                   `_@�>����?-            @T@              #                 ����? =[y��?&             Q@                                  �?�L���?            �B@        ������������������������       �                     $@                                   �?�����H�?             ;@        ������������������������       �                     .@                                  �Y@      �?             (@       ������������������������       �                     @               "                    \@���Q��?             @               !                    @O@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ?@        %       &                    ^@�θ�?             *@        ������������������������       �                      @        '       (                    �?�C��2(�?             &@        ������������������������       �                     @        )       *                    `@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        -       2                    �?"pc�
�?             &@       .       /                     Q@�<ݚ�?             "@        ������������������������       �                     @        0       1                    �Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        6       C                 pff�?���!pc�?.            @S@       7       B                    �?@4և���?"             L@        8       =                    �?�	j*D�?	             *@       9       :                    �?և���X�?             @        ������������������������       �                      @        ;       <                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        >       ?                     M@r�q��?             @        ������������������������       �                     @        @       A                   `Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �E@        D       G                    �K@��s����?             5@        E       F                    `@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        I       �                    �?�;����?�            �x@        J       {       
             �?b��H���?a            �b@       K       v                   �a@�����?K            �\@       L       m       	             �?|�|k6��?7            �U@       M       N                   �U@�̚��?(            �N@        ������������������������       �                     @        O       b                    @M@P̏����?'            �L@       P       W                    �?�p ��?            �D@        Q       V                   �q@      �?              @       R       U                 ����?z�G�z�?             @       S       T                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        X       _                    �?�FVQ&�?            �@@       Y       ^                    �E@�g�y��?             ?@       Z       ]                    �?��S�ۿ?             .@       [       \                   �r@�C��2(�?	             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        `       a                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        c       f                    @O@      �?
             0@        d       e                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        g       l                   �\@�<ݚ�?             "@        h       k                   �c@���Q��?             @       i       j                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        n       o                   �\@$��m��?             :@        ������������������������       �                     @        p       s                    @L@��s����?             5@       q       r                    @�IєX�?
             1@       ������������������������       �        	             0@        ������������������������       �                     �?        t       u                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        w       x                    �? 7���B�?             ;@       ������������������������       �                     8@        y       z                   p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        |       }                   `\@�ʻ����?             A@        ������������������������       �                     @        ~                            H@���@M^�?             ?@        ������������������������       �                     @        �       �                    �?      �?             8@       �       �                    �?      �?             (@       ������������������������       �                     @        �       �                 ����?���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    b@      �?             (@       �       �                   �b@�����H�?             "@        �       �                     L@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �L@ĭ����?�            @o@       �       �                   @g@�q-�?z             j@       �       �                   �O@��ɶ�"�?y            �i@        �       �                   �Z@�q�q�?             @        ������������������������       �                      @        �       �                 ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�����?v             i@       �       �       	             �?�=
ףp�?Z             d@        �       �                   @[@ ����?&            @P@        �       �       
             �?z�G�z�?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   @Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        "             N@        ������������������������       �        4            �W@        �       �                 433�?� ��1�?            �D@       �       �                    �?(N:!���?            �A@       �       �                    \@؇���X�?             <@        �       �                     H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   d@HP�s��?             9@        ������������������������       �                     *@        �       �                   p@r�q��?             (@        �       �                    �?      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                     I@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@����X�?!             E@        �       �                   �?�\��N��?             3@       �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �                   �c@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   Pc@      �?              @        �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?���}<S�?             7@       �       �                   �j@���7�?             6@        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B  �%փmM�?+�>IY�?��y��y�?�a�a�?�{�ո�?��P��?l(�����?(������?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?DDDDDD�?��?�`��`��?ysB�n�?��k���?              �?qBJ�eD�?�[���?�������?ffffff�?h/�����?�Kh/��?�������?�������?L�Ϻ��?}���g�?              �?�q�q�?�q�q�?              �?      �?      �?              �?333333�?�������?      �?      �?              �?      �?              �?                      �?�؉�؉�?ى�؉��?      �?        F]t�E�?]t�E�?              �?�������?�������?      �?                      �?              �?F]t�E�?/�袋.�?�q�q�?9��8���?              �?      �?      �?      �?                      �?              �?      �?              �?        F]t�E�?t�E]t�?n۶m۶�?�$I�$I�?vb'vb'�?;�;��?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �a�a�?z��y���?�$I�$I�?۶m۶m�?              �?      �?                      �? �'�n�?�=�ѻ"�?�|����?�����?^Cy�5�?Q^Cy��?;���C��?�2)^ �?�u�y���??�%C���?      �?        ��Gp�??���#�?��+Q��?Q��+Q�?      �?      �?�������?�������?      �?      �?      �?                      �?      �?                      �?|���?>����?�B!��?��{���?�?�������?F]t�E�?]t�E�?              �?      �?                      �?              �?      �?      �?              �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?                      �?�q�q�?9��8���?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�N��N��?vb'vb'�?              �?z��y���?�a�a�?�?�?      �?                      �?      �?      �?              �?      �?        h/�����?	�%����?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?<<<<<<�?              �?�s�9��?�c�1��?      �?              �?      �?      �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        y�&1��?9��v���?��؉���?�;�;�?�pK͆��?�{����?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?g��1��?���@��?�������?������y? �����? �����?�������?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ������?������?|�W|�W�?�A�A�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?        q=
ףp�?{�G�z�?      �?        �������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?�m۶m��?�$I�$I�?�5��P�?y�5���?F]t�E�?t�E]t�?      �?              �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?ӛ���7�?d!Y�B�?�.�袋�?F]t�E�?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJcʚhG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B@5         �                    �?&I,|-��?�           ��@              w       	             �?�h�C�J�?           �y@              ^                   �b@�G�2��?�            �w@              G       
             �?p`�i0�?�            �s@              *                 ����?���x���?�            �p@                                   �?����?H             ]@                                  @M@,sI�v�?9            �V@                                  �?&y�X���?#             M@       	                          �s@      �?             F@       
                        ����?d}h���?             E@        ������������������������       �        	             (@                                   �?�z�G��?             >@                                  �?�X����?             6@        ������������������������       �                     @                                  �`@r�q��?	             2@       ������������������������       �                     (@                                  �Z@      �?             @        ������������������������       �                      @                                   b@      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             ,@        ������������������������       �                     @@                                  �i@�	j*D�?             :@       ������������������������       �                     (@                )                    b@և���X�?             ,@       !       $                   �_@���!pc�?             &@        "       #                    ]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        %       (                   �k@؇���X�?             @        &       '                   �j@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        +       ,                    �?��F��?i            `c@        ������������������������       �                     @@        -       :                    �?@;�"�?W            �^@        .       /                    �?\-��p�?             =@        ������������������������       �        	             ,@        0       5                    �?������?             .@       1       2                   @a@z�G�z�?             $@       ������������������������       �                     @        3       4                    Y@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        6       7                 `ff�?���Q��?             @        ������������������������       �                      @        8       9                   @p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ;       D                   @b@`�q�0ܴ?C            �W@       <       C                    \@hl �&�?A             W@        =       >                    �?��a�n`�?             ?@       ������������������������       �                     6@        ?       @                   �[@�q�q�?             "@       ������������������������       �                     @        A       B                     M@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        ,            �N@        E       F                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        H       M                    �?t/*�?$            �G@        I       J                 ����?      �?              @        ������������������������       �                     @        K       L                    o@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        N       O                    `@��-�=��?            �C@        ������������������������       �        
             0@        P       ]                   �r@�㙢�c�?             7@       Q       X                   �`@��2(&�?             6@       R       W                    �?      �?             0@        S       T                    �Q@z�G�z�?             @        ������������������������       �                     @        U       V                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@        Y       Z                    �?�q�q�?             @        ������������������������       �                     @        [       \                 ���@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                   �g@�q�q�?"             N@        ������������������������       �                     0@        a       p                   �o@�eP*L��?             F@       b       k                    `@�	j*D�?             :@       c       d       
             �?�q�q�?	             (@        ������������������������       �                     @        e       f                    �?����X�?             @        ������������������������       �                      @        g       h                     I@���Q��?             @        ������������������������       �                      @        i       j                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        l       o                 ����?@4և���?             ,@        m       n                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        q       v       
             �?�����H�?
             2@       r       s                   �r@�IєX�?	             1@       ������������������������       �                     (@        t       u                   @^@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        x                          �b@���|���?            �@@       y       z                   �[@      �?             <@        ������������������������       �                     @        {       |                   �\@�J�4�?             9@        ������������������������       �                     @        }       ~                    @���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��+Q���?�            0t@       �       �                   h@l�b�G��?�            �l@       �       �                   @[@ (��?�            @l@        �       �                    �F@@�0�!��?             1@       ������������������������       �                     (@        �       �                    c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       	             �?�}�+r��?�             j@        �       �                   �a@�8��8��?<             X@        �       �                    �?�(\����?             D@       ������������������������       �                     B@        �       �                    �?      �?             @       �       �                    @L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �t@      �?%             L@       �       �                 ���@$�q-�?#             J@       �       �                    �?@�E�x�?             �H@       ������������������������       �                     F@        �       �                   0i@z�G�z�?             @        ������������������������       �                     @        �       �                 033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? T���v�?L            @\@       �       �                    �?�|1)�?G            �Z@       �       �                   �? f^8���?E            �Y@       ������������������������       �        ;            @U@        �       �                 pff�?r�q��?
             2@        �       �                   p`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @P@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?d��4�o�?:            �W@       �       �                    �?�	j*D�?/            �S@       �       �                 @33�?��$�4��?$            �M@       �       �                   �`@t��ճC�?             F@        ������������������������       �                     5@        �       �                    �?�LQ�1	�?             7@       �       �                   pf@      �?
             0@       �       �                   �c@��S�ۿ?	             .@       ������������������������       �                     &@        �       �                   0i@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    T@؇���X�?             @        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �d@�q�q�?	             .@       �       �                   �j@r�q��?             (@       �       �                 ����?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    k@D�n�3�?             3@        ������������������������       �                     @        �       �                    �D@և���X�?             ,@        ������������������������       �                     @        �       �                    �L@���!pc�?             &@       ������������������������       �                     @        �       �                   f@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   `\@������?             1@       ������������������������       �                     (@        �       �                   0c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�BP  �"z?+�?���B`��?ؿ$J��?
�6x-�?�)��ԟ�?���
X�?J�-�?��6b]z�?Q�Ѿj��?6�%����?�rO#,��?O#,�4��?��I��I�?l�l��?�i��F�?��FX��?      �?      �?۶m۶m�?I�$I�$�?              �?333333�?ffffff�?]t�E]�?�E]t��?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?                      �?              �?;�;��?vb'vb'�?              �?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?mЦm�?Y���/Y�?              �?�h
���?����/��?�{a���?a����?              �?�?wwwwww�?�������?�������?              �?�������?333333�?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        W�+�ɥ?��F}g��?Y�B��?ozӛ���?�c�1Ƹ?�s�9��?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?W�+���?�;����?      �?      �?              �?�������?�������?      �?                      �?�A�A�?}˷|˷�?              �?d!Y�B�?�7��Mo�?t�E]t�?��.���?      �?      �?�������?�������?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?vb'vb'�?;�;��?�������?�������?              �?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?        �q�q�?�q�q�?�?�?              �?�������?�������?      �?                      �?      �?        ]t�E]�?F]t�E�?      �?      �?              �?�z�G��?{�G�z�?              �?�.�袋�?F]t�E�?      �?                      �?              �?9�FͿ�?_��� �?�Gp��?p�}��?H���?x�!���?ZZZZZZ�?�������?      �?        �������?333333�?              �?      �?        �5��P�?(�����?UUUUUU�?UUUUUU�?333333�?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�؉�؉�?;�;��?և���X�?9/���?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?      �?      �?      �?                      �?6h�e�&�?4��A�/�?W�9�&�?"5�x+��?H%�e�?��VCӝ?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �������?�?      �?                      �?      �?              �?                      �?�8�{n��?Ҏ#��?vb'vb'�?;�;��?#h8����?u_[4�?�E]t��?t�E]t�?      �?        ��Moz��?Y�B��?      �?      �?�������?�?      �?              �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?�q�q�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        (������?l(�����?              �?�$I�$I�?۶m۶m�?              �?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?        �?xxxxxx�?              �?�������?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5&]hG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKㅔh��B�8         �                    �?"�\�&U�?�           ��@              )                    �?ʋ�A��?           pz@               $                   �c@և���X�?)            �O@                                  �?���|���?#            �K@                                  0c@և���X�?             <@                                 `X@      �?             4@        ������������������������       �                      @                      	             �?r�q��?             2@       	       
                   �`@      �?             (@        ������������������������       �                      @                                    P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �N@      �?              @       ������������������������       �                     @                                ���@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  h@PN��T'�?             ;@                                  �V@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                   �?���}<S�?             7@                               ����?�X�<ݺ?             2@                                   �H@؇���X�?             @                                  @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@                #                   @_@z�G�z�?             @       !       "                   hs@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        %       &                    �?      �?              @        ������������������������       �                     @        '       (                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        *       e                    �?���Hx�?�            �v@        +       :                   �a@t/*�?Y            �a@       ,       -                   �]@xdQ�m��?1            @T@       ������������������������       �                     H@        .       1                    �?6YE�t�?            �@@        /       0                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        2       9                    �? 7���B�?             ;@       3       8                    �?�X�<ݺ?             2@        4       7                    �?z�G�z�?             @        5       6       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     "@        ;       V                   a@^n����?(             N@       <       =                   `\@H�z�G�?             D@        ������������������������       �                     "@        >       ?                   �]@`՟�G��?             ?@        ������������������������       �                      @        @       Q                    �?l��[B��?             =@       A       N       
             �?\X��t�?             7@       B       G                    �?��.k���?             1@       C       F                   �`@���Q��?             $@       D       E                    p@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        H       I                    �?����X�?             @        ������������������������       �                      @        J       K                   @]@���Q��?             @        ������������������������       �                      @        L       M                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        O       P                   �_@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        R       S                   @_@�q�q�?             @        ������������������������       �                     �?        T       U                    �L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        W       ^                    �?ףp=
�?             4@       X       ]                   �a@$�q-�?	             *@       Y       \                   �j@r�q��?             @        Z       [       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        _       d                    �?؇���X�?             @       `       a                   @c@z�G�z�?             @        ������������������������       �                      @        b       c                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        f       �                    �R@h�j��l�?�            `k@       g       �                    �? '��h�?�            @k@       h       �                   pb@ ��Ou��?b            �c@       i       n                    �?�2c�$��?[             b@        j       m                   P`@XB���?             =@        k       l                   �\@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        o       x                    \@�8���?F             ]@        p       w                    �?�q�q�?             (@       q       v                    �?z�G�z�?             $@       r       s                    �I@���Q��?             @        ������������������������       �                      @        t       u                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        y       �                    �? pƵHP�??             Z@       z       �                    �?`��>�ϗ?2            @U@       {       |                   Xp@`׀�:M�?+            �R@       ������������������������       �                     C@        }       �                 ����?������?             B@        ~                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        ������������������������       �                     &@        �       �                   �_@�}�+r��?             3@        �       �                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                   �Z@���!pc�?             &@        ������������������������       �                      @        �       �                    q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        (             O@        ������������������������       �                     �?        �       �                   @E@Σq���?�            ps@        �       �                     O@     ��?             @@       �       �                    �?�LQ�1	�?             7@        �       �                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�}�+r��?             3@       ������������������������       �                     &@        �       �                 `ff�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ����?X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �]@�q�q�?             @        ������������������������       �                      @        �       �                     Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?īr4e�?�            pq@       �       �                   �X@`� x��?�            �l@        ������������������������       �                     �?        �       �       
             �?�`z����?�            `l@       �       �                    �?�8��8��?m             e@       �       �       	             �?`�߻�ɒ?H             [@        ������������������������       �                      @        �       �                    @L@ �ׁsF�?A             Y@       ������������������������       �        :             W@        �       �                   �?      �?              @       ������������������������       �                     @        �       �                 pff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 033�?d��0u��?%             N@       �       �                   �b@Hm_!'1�?            �H@       �       �                     N@`�q�0ܴ?            �G@       �       �                    �? ���J��?            �C@       �       �                    �? 7���B�?             ;@        ������������������������       �                      @        �       �                   �n@`2U0*��?             9@       ������������������������       �                     5@        �       �                    �H@      �?             @        ������������������������       �                      @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?���#�İ?&            �M@       �       �                     O@h�����?#             L@       ������������������������       �        !             J@        �       �                    a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @�q�q�?             �I@       �       �                 ����?`�Q��?             I@       �       �       	             �?�LQ�1	�?             G@       �       �                    �?*O���?             B@       ������������������������       �                     0@        �       �                    �?��Q��?             4@       �       �                   `\@     ��?             0@       �       �                    @I@���!pc�?             &@       ������������������������       �                     @        �       �                    �N@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   d@z�G�z�?             @        ������������������������       �                      @        �       �                   �e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    d@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hi�B0  ��j��`�?:�J;�O�?�1�����?�s�HO�?۶m۶m�?�$I�$I�?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?      �?              �?�������?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?h/�����?&���^B�?      �?      �?              �?      �?        d!Y�B�?ӛ���7�?�q�q�?��8��8�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?�������?�������?      �?      �?      �?                      �?              �?      �?      �?      �?        �������?�������?              �?      �?        9��8��?9��8���?W�+���?�;����?X�<ݚ�?�5?,R�?              �?e�M6�d�?'�l��&�?UUUUUU�?UUUUUU�?              �?      �?        h/�����?	�%����?�q�q�?��8��8�?�������?�������?      �?      �?      �?                      �?              �?              �?              �?DDDDDD�?�������?333333�?ffffff�?              �?�1�c��?�s�9��?      �?        ���=��?GX�i���?!Y�B�?��Moz��?�?�������?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?�m۶m��?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?        �������?�������?;�;��?�؉�؉�?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?x��m���?H�!��d�?�w� z|�?���]8��?�i�i�?.��-���?�y�!���?cH�-�t�?�{a���?GX�i���?      �?      �?              �?      �?                      �?a���{�?j��FX�?UUUUUU�?UUUUUU�?�������?�������?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ;�;��?'vb'vb�?�?�������?к����?��L��?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?              �?(�����?�5��P�?UUUUUU�?UUUUUU�?              �?      �?                      �?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?                      �?      �?        !�J���?|_��oH�?      �?      �?Y�B��?��Moz��?      �?      �?      �?                      �?(�����?�5��P�?              �?      �?      �?              �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�f���?��|Hw2�?�YLg1��?g1��t�?              �?�s���?��gG�?UUUUUU�?UUUUUU�?B{	�%��?h/�����?      �?        �G�z��?{�G�z�?      �?              �?      �?      �?              �?      �?              �?      �?        �?�������?Y�Cc�?9/���?��F}g��?W�+�ɥ?��-��-�?�A�A�?	�%����?h/�����?      �?        ���Q��?{�G�z�?      �?              �?      �?      �?              �?      �?      �?                      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?/�袋.�?      �?                      �?��N��?'u_[�?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?��(\���?{�G�z�?Nozӛ��?d!Y�B�?�q�q�?�q�q�?      �?        ffffff�?�������?      �?      �?t�E]t�?F]t�E�?              �?333333�?�������?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?333333�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�K6ShG        hNhG        hNhMKhOKhPh)h,K ��h.��R�(KK��hi�C              �?�t�bh\hnhWC       ���R�hrKhshvKh)h,K ��h.��R�(KK��hW�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��B�;         �                    �?4�5����?�           ��@              �       	             �?@�B��q�?           @{@              ^                   �`@.�P*�b�?�            y@               %                    �?@�҇��?z            �g@               
                 ����?X�Emq�?!            �J@               	                    �?@4և���?             ,@                                  �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �Q@��Zy�?            �C@                                  �c@      �?             (@       ������������������������       �                      @                                  �d@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                  `\@l��
I��?             ;@                                033@և���X�?             @                                 @a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                   �?z�G�z�?             4@        ������������������������       �                     @               "                    �?������?             1@              !                    �?$�q-�?	             *@                                  �?      �?              @        ������������������������       �                     @                                  �k@z�G�z�?             @        ������������������������       �                      @                                   Pm@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        #       $                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        &       3                    �?Xș���?Y            �`@        '       2                    �?      �?             0@       (       1                    �?�n_Y�K�?	             *@       )       *                    �?z�G�z�?             $@        ������������������������       �                     @        +       ,                 ����?�q�q�?             @        ������������������������       �                     @        -       .                 ����?�q�q�?             @        ������������������������       �                     �?        /       0                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        4       ;                    @J@��5Վ3�?N            �]@        5       :                    �? �q�q�?             H@        6       7                   �`@z�G�z�?             $@       ������������������������       �                     @        8       9                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     C@        <       E                   @X@O�o9%�?/            �Q@        =       >                   �Y@      �?              @        ������������������������       �                     �?        ?       @                   @_@����X�?             @        ������������������������       �                     �?        A       B                   l@r�q��?             @        ������������������������       �                     @        C       D                    T@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        F       Y                    �?�? Da�?*            �O@       G       X                    �?�:�]��?#            �I@       H       S                    @(N:!���?            �A@       I       J                    �?��S�ۿ?             >@        ������������������������       �                     &@        K       L                 433�?�KM�]�?             3@        ������������������������       �                     �?        M       R                    �?�X�<ݺ?             2@       N       Q                 `ff�?$�q-�?             *@        O       P                 ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        T       W                   �_@���Q��?             @       U       V                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        Z       ]                   �[@�q�q�?             (@       [       \                    @L@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        _       v                    �?��Hw��?�            �j@       `       e                    �?��j��Ѳ?`            �c@        a       d                    �R@�r����?             .@       b       c                    �?@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        f       u                    �R@�J�T�?X            �a@       g       t                 ����?`����֜?W            �a@        h       i                   a@h㱪��?"            �K@       ������������������������       �                    �A@        j       o                    �?ףp=
�?             4@       k       n                    �?�C��2(�?             &@       l       m                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        p       q                   @b@�����H�?             "@        ������������������������       �                     @        r       s                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        5            @U@        ������������������������       �                      @        w       �                    �?4և����?!             L@        x       �       
             �?� �	��?             9@       y       z                    �?�q�q�?             5@        ������������������������       �                      @        {       �                    �?p�ݯ��?             3@        |       }                   c@X�<ݚ�?             "@        ������������������������       �                     @        ~                          �c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �b@`Jj��?             ?@       ������������������������       �                     =@        ������������������������       �                      @        �       �                   �`@<=�,S��?            �A@       �       �                    �B@      �?             <@        ������������������������       �                     �?        �       �                   �Z@�<ݚ�?             ;@        ������������������������       �                     @        �       �                    �?      �?             8@        �       �                 033�?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?P���Q�?	             4@       ������������������������       �                     ,@        �       �                    @L@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        �       �                   s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @L@��H�&p�?�            �r@       �       �                    �?��x��?�            @i@       �       �       	             �?���.�6�?|             g@       �       �       
             �?�����?I            @Z@        �       �                    �?>a�����?$            �I@       �       �                   @E@���H��?             E@        �       �                   @_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   pj@�}�+r��?             C@        ������������������������       �        	             0@        �       �                    �?�C��2(�?             6@       �       �                    �?���N8�?             5@        ������������������������       �                      @        �       �                   �j@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        �       �                    @F@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                     G@ 7���B�?%             K@        ������������������������       �                     9@        �       �                    �? 	��p�?             =@       �       �                    �?$�q-�?             :@       �       �                   @[@���}<S�?             7@        ������������������������       �                     �?        �       �                 ����?���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �g@pY���D�?3            �S@       ������������������������       �        1            �R@        �       �                    �D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �E@b�2�tk�?             2@        ������������������������       �                      @        �       �                    �?     ��?             0@       �       �                   `]@r�q��?             (@        ������������������������       �                     �?        �       �                   `@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   d@     ��?9             X@        �       �                   `@�θ�?             *@        ������������������������       �                     @        �       �                   `_@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �c@�0���?1            �T@       �       �                   �o@�+$�jP�?             K@       �       �       
             �?�g�y��?             ?@       �       �                 ����?�nkK�?             7@       ������������������������       �                     4@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0q@�û��|�?             7@        �       �                   Hp@�����H�?             "@        �       �                    p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Z@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?П[;U��?             =@        ������������������������       �                     $@        �       �       
             �?�����?             3@       �       �                   `d@r�q��?             (@       ������������������������       �                      @        �       �                   0e@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    e@և���X�?             @        ������������������������       �                     @        �       �                   �h@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�b�'      h�h)h,K ��h.��R�(KK�KK��hi�B�   Np	�?���Gw{�?��[����?���[��?��*m���?�N����?}g���Q�?!&W�+�?�}�	��?5�x+��?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?� � �?\��[���?      �?      �?              �?      �?      �?      �?                      �?Lh/����?h/�����?۶m۶m�?�$I�$I�?333333�?�������?              �?      �?                      �?�������?�������?      �?        xxxxxx�?�?�؉�؉�?;�;��?      �?      �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        �\y@���?Ũ�oS��?      �?      �?;�;��?ى�؉��?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?�k"�k"�?e�e��?UUUUUU�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?��RO�o�?�D+l$�?      �?      �?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?AA�?�������?�?}}}}}}�?�A�A�?|�W|�W�?�?�������?              �?(�����?�k(���?      �?        �q�q�?��8��8�?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?�q�q�?r�q��?      �?                      �?              �?0x,�ն?��pB%�?A����?|DN���?�?�������?�$I�$I�?n۶m۶�?      �?                      �?      �?        ��V؜?(�K=�?�A�A�?�������?��)A��?־a���?              �?�������?�������?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        n۶m۶�?%I�$I��?)\���(�?�Q����?UUUUUU�?UUUUUU�?              �?Cy�5��?^Cy�5�?�q�q�?r�q��?              �?�������?�������?      �?                      �?333333�?ffffff�?      �?                      �?      �?        �B!��?���{��?              �?      �?        �A�A�?X|�W|��?      �?      �?              �?9��8���?�q�q�?              �?      �?      �?      �?      �?      �?                      �?ffffff�?�������?      �?        �������?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?��o�j�?�IA��U�?�S� w��?�be�F�?���7���?Y�B��?=��<���?�a�a�?�������?�?�0�0�?��y��y�?      �?      �?              �?      �?        �5��P�?(�����?      �?        ]t�E�?F]t�E�?��y��y�?�a�a�?      �?        �5��P�?(�����?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        	�%����?h/�����?      �?        ������?�{a���?�؉�؉�?;�;��?ӛ���7�?d!Y�B�?              �?�.�袋�?F]t�E�?      �?                      �?      �?              �?        a~W��0�?�3���?      �?        333333�?�������?      �?                      �?�8��8��?9��8���?              �?      �?      �?�������?UUUUUU�?              �?]t�E�?F]t�E�?              �?      �?              �?      �?      �?                      �?      �?      �?�؉�؉�?ى�؉��?              �?۶m۶m�?�$I�$I�?              �?      �?        o4u~�!�?"�%��?/�����?B{	�%��?��{���?�B!��?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        8��Moz�?��,d!�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?n۶m۶�?�$I�$I�?              �?      �?        �{a���?��=���?      �?        ^Cy�5�?Q^Cy��?UUUUUU�?�������?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?�t�bubhhubehhub.